library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0fcc287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49c0fcc2",
    18 => x"48d8e3c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"d8e3c287",
    25 => x"d4e3c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e8c187f7",
    29 => x"e3c287fb",
    30 => x"e3c24dd8",
    31 => x"ad744cd8",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"8148731e",
    65 => x"c502a973",
    66 => x"05531287",
    67 => x"4f2687f6",
    68 => x"711e731e",
    69 => x"4b66c84a",
    70 => x"718bc149",
    71 => x"87cf0299",
    72 => x"d4ff4812",
    73 => x"49737808",
    74 => x"99718bc1",
    75 => x"2687f105",
    76 => x"0e4f264b",
    77 => x"0e5c5b5e",
    78 => x"d4ff4a71",
    79 => x"4b66cc4c",
    80 => x"718bc149",
    81 => x"87ce0299",
    82 => x"6c7cffc3",
    83 => x"c1497352",
    84 => x"0599718b",
    85 => x"4c2687f2",
    86 => x"4f264b26",
    87 => x"ff1e731e",
    88 => x"ffc34bd4",
    89 => x"c34a6b7b",
    90 => x"496b7bff",
    91 => x"b17232c8",
    92 => x"6b7bffc3",
    93 => x"7131c84a",
    94 => x"7bffc3b2",
    95 => x"32c8496b",
    96 => x"4871b172",
    97 => x"4f264b26",
    98 => x"5c5b5e0e",
    99 => x"4d710e5d",
   100 => x"754cd4ff",
   101 => x"98ffc348",
   102 => x"e3c27c70",
   103 => x"c805bfd8",
   104 => x"4866d087",
   105 => x"a6d430c9",
   106 => x"4966d058",
   107 => x"487129d8",
   108 => x"7098ffc3",
   109 => x"4966d07c",
   110 => x"487129d0",
   111 => x"7098ffc3",
   112 => x"4966d07c",
   113 => x"487129c8",
   114 => x"7098ffc3",
   115 => x"4866d07c",
   116 => x"7098ffc3",
   117 => x"d049757c",
   118 => x"c3487129",
   119 => x"7c7098ff",
   120 => x"f0c94b6c",
   121 => x"ffc34aff",
   122 => x"87cf05ab",
   123 => x"6c7c7149",
   124 => x"028ac14b",
   125 => x"ab7187c5",
   126 => x"7387f202",
   127 => x"264d2648",
   128 => x"264b264c",
   129 => x"49c01e4f",
   130 => x"c348d4ff",
   131 => x"81c178ff",
   132 => x"a9b7c8c3",
   133 => x"2687f104",
   134 => x"5b5e0e4f",
   135 => x"c00e5d5c",
   136 => x"f7c1f0ff",
   137 => x"c0c0c14d",
   138 => x"4bc0c0c0",
   139 => x"c487d6ff",
   140 => x"c04cdff8",
   141 => x"fd49751e",
   142 => x"86c487ce",
   143 => x"c005a8c1",
   144 => x"d4ff87e5",
   145 => x"78ffc348",
   146 => x"e1c01e73",
   147 => x"49e9c1f0",
   148 => x"c487f5fc",
   149 => x"05987086",
   150 => x"d4ff87ca",
   151 => x"78ffc348",
   152 => x"87cb48c1",
   153 => x"c187defe",
   154 => x"c6ff058c",
   155 => x"2648c087",
   156 => x"264c264d",
   157 => x"0e4f264b",
   158 => x"0e5c5b5e",
   159 => x"c1f0ffc0",
   160 => x"d4ff4cc1",
   161 => x"78ffc348",
   162 => x"f849fcca",
   163 => x"4bd387d9",
   164 => x"49741ec0",
   165 => x"c487f1fb",
   166 => x"05987086",
   167 => x"d4ff87ca",
   168 => x"78ffc348",
   169 => x"87cb48c1",
   170 => x"c187dafd",
   171 => x"dfff058b",
   172 => x"2648c087",
   173 => x"264b264c",
   174 => x"0000004f",
   175 => x"00444d43",
   176 => x"43484453",
   177 => x"69616620",
   178 => x"000a216c",
   179 => x"52524549",
   180 => x"00000000",
   181 => x"00495053",
   182 => x"74697257",
   183 => x"61662065",
   184 => x"64656c69",
   185 => x"5e0e000a",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"d0fc4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"c7fa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087ecfd",
   195 => x"87e8c148",
   196 => x"7087c9f9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fd87c802",
   200 => x"48c087d5",
   201 => x"7587d1c1",
   202 => x"4cf1c07b",
   203 => x"7087eafb",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87c8f949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"db48c187",
   215 => x"d748c087",
   216 => x"05acc287",
   217 => x"c0cb87ca",
   218 => x"87fbf449",
   219 => x"87c848c0",
   220 => x"fe058cc1",
   221 => x"48c087f6",
   222 => x"4c264d26",
   223 => x"4f264b26",
   224 => x"5c5b5e0e",
   225 => x"d0ff0e5d",
   226 => x"d0e5c04d",
   227 => x"c24cc0c1",
   228 => x"c148d8e3",
   229 => x"49d4cb78",
   230 => x"c787ccf4",
   231 => x"f97dc24b",
   232 => x"7dc387e3",
   233 => x"49741ec0",
   234 => x"c487ddf7",
   235 => x"05a8c186",
   236 => x"c24b87c1",
   237 => x"87cb05ab",
   238 => x"f349cccb",
   239 => x"48c087e9",
   240 => x"c187f6c0",
   241 => x"d4ff058b",
   242 => x"87dafc87",
   243 => x"58dce3c2",
   244 => x"cd059870",
   245 => x"c01ec187",
   246 => x"d0c1f0ff",
   247 => x"87e8f649",
   248 => x"d4ff86c4",
   249 => x"78ffc348",
   250 => x"c287eec4",
   251 => x"c258e0e3",
   252 => x"48d4ff7d",
   253 => x"c178ffc3",
   254 => x"264d2648",
   255 => x"264b264c",
   256 => x"5b5e0e4f",
   257 => x"710e5d5c",
   258 => x"4cffc34d",
   259 => x"744bd4ff",
   260 => x"48d0ff7b",
   261 => x"7478c3c4",
   262 => x"c01e757b",
   263 => x"d8c1f0ff",
   264 => x"87e4f549",
   265 => x"987086c4",
   266 => x"cb87cb02",
   267 => x"f6f149d8",
   268 => x"c048c187",
   269 => x"7b7487ee",
   270 => x"c87bfec3",
   271 => x"66d41ec0",
   272 => x"87ccf349",
   273 => x"7b7486c4",
   274 => x"7b747b74",
   275 => x"4ae0dad8",
   276 => x"056b7b74",
   277 => x"8ac187c5",
   278 => x"7487f505",
   279 => x"48d0ff7b",
   280 => x"48c078c2",
   281 => x"4c264d26",
   282 => x"4f264b26",
   283 => x"5c5b5e0e",
   284 => x"86fc0e5d",
   285 => x"d4ff4b71",
   286 => x"c57ec04c",
   287 => x"4adfcdee",
   288 => x"6c7cffc3",
   289 => x"a8fec348",
   290 => x"87f8c005",
   291 => x"9b734d74",
   292 => x"d487cc02",
   293 => x"49731e66",
   294 => x"c487d8f2",
   295 => x"ff87d486",
   296 => x"d1c448d0",
   297 => x"4a66d478",
   298 => x"c17dffc3",
   299 => x"87f8058a",
   300 => x"c35aa6d8",
   301 => x"737c7cff",
   302 => x"87c5059b",
   303 => x"d048d0ff",
   304 => x"7e4ac178",
   305 => x"fe058ac1",
   306 => x"486e87f6",
   307 => x"4d268efc",
   308 => x"4b264c26",
   309 => x"731e4f26",
   310 => x"c04a711e",
   311 => x"48d4ff4b",
   312 => x"ff78ffc3",
   313 => x"c3c448d0",
   314 => x"48d4ff78",
   315 => x"7278ffc3",
   316 => x"f0ffc01e",
   317 => x"f249d1c1",
   318 => x"86c487ce",
   319 => x"d2059870",
   320 => x"1ec0c887",
   321 => x"fd4966cc",
   322 => x"86c487e2",
   323 => x"d0ff4b70",
   324 => x"7378c248",
   325 => x"264b2648",
   326 => x"5b5e0e4f",
   327 => x"c00e5d5c",
   328 => x"f0ffc01e",
   329 => x"f149c9c1",
   330 => x"1ed287de",
   331 => x"49e8e3c2",
   332 => x"c887f9fc",
   333 => x"c14cc086",
   334 => x"acb7d284",
   335 => x"c287f804",
   336 => x"bf97e8e3",
   337 => x"99c0c349",
   338 => x"05a9c0c1",
   339 => x"c287e7c0",
   340 => x"bf97efe3",
   341 => x"c231d049",
   342 => x"bf97f0e3",
   343 => x"7232c84a",
   344 => x"f1e3c2b1",
   345 => x"b14abf97",
   346 => x"ffcf4c71",
   347 => x"c19cffff",
   348 => x"c134ca84",
   349 => x"e3c287e7",
   350 => x"49bf97f1",
   351 => x"99c631c1",
   352 => x"97f2e3c2",
   353 => x"b7c74abf",
   354 => x"c2b1722a",
   355 => x"bf97ede3",
   356 => x"9dcf4d4a",
   357 => x"97eee3c2",
   358 => x"9ac34abf",
   359 => x"e3c232ca",
   360 => x"4bbf97ef",
   361 => x"b27333c2",
   362 => x"97f0e3c2",
   363 => x"c0c34bbf",
   364 => x"2bb7c69b",
   365 => x"81c2b273",
   366 => x"307148c1",
   367 => x"48c14970",
   368 => x"4d703075",
   369 => x"84c14c72",
   370 => x"c0c89471",
   371 => x"cc06adb7",
   372 => x"b734c187",
   373 => x"b7c0c82d",
   374 => x"f4ff01ad",
   375 => x"26487487",
   376 => x"264c264d",
   377 => x"0e4f264b",
   378 => x"5d5c5b5e",
   379 => x"c286fc0e",
   380 => x"c048d0ec",
   381 => x"c8e4c278",
   382 => x"fb49c01e",
   383 => x"86c487d8",
   384 => x"c5059870",
   385 => x"c948c087",
   386 => x"4dc087d2",
   387 => x"48ccf1c2",
   388 => x"e4c278c1",
   389 => x"e1c04afe",
   390 => x"4bc849f4",
   391 => x"7087c7eb",
   392 => x"87c60598",
   393 => x"48ccf1c2",
   394 => x"e5c278c0",
   395 => x"e2c04ada",
   396 => x"4bc849c0",
   397 => x"7087efea",
   398 => x"87c60598",
   399 => x"48ccf1c2",
   400 => x"f1c278c0",
   401 => x"c002bfcc",
   402 => x"ebc287fd",
   403 => x"c24dbfce",
   404 => x"bf9fc6ec",
   405 => x"d6c5487e",
   406 => x"c705a8ea",
   407 => x"ceebc287",
   408 => x"87ce4dbf",
   409 => x"e9ca486e",
   410 => x"c502a8d5",
   411 => x"c748c087",
   412 => x"e4c287ea",
   413 => x"49751ec8",
   414 => x"c487dbf9",
   415 => x"05987086",
   416 => x"48c087c5",
   417 => x"c287d5c7",
   418 => x"c04adae5",
   419 => x"c849cce2",
   420 => x"87d2e94b",
   421 => x"c8059870",
   422 => x"d0ecc287",
   423 => x"d878c148",
   424 => x"fee4c287",
   425 => x"d8e2c04a",
   426 => x"e84bc849",
   427 => x"987087f8",
   428 => x"87c5c002",
   429 => x"e3c648c0",
   430 => x"c6ecc287",
   431 => x"c149bf97",
   432 => x"c005a9d5",
   433 => x"ecc287cd",
   434 => x"49bf97c7",
   435 => x"02a9eac2",
   436 => x"c087c5c0",
   437 => x"87c4c648",
   438 => x"97c8e4c2",
   439 => x"c3487ebf",
   440 => x"c002a8e9",
   441 => x"486e87ce",
   442 => x"02a8ebc3",
   443 => x"c087c5c0",
   444 => x"87e8c548",
   445 => x"97d3e4c2",
   446 => x"059949bf",
   447 => x"c287ccc0",
   448 => x"bf97d4e4",
   449 => x"02a9c249",
   450 => x"c087c5c0",
   451 => x"87ccc548",
   452 => x"97d5e4c2",
   453 => x"ecc248bf",
   454 => x"4c7058cc",
   455 => x"c288c148",
   456 => x"c258d0ec",
   457 => x"bf97d6e4",
   458 => x"c2817549",
   459 => x"bf97d7e4",
   460 => x"7232c84a",
   461 => x"f0c27ea1",
   462 => x"786e48e8",
   463 => x"97d8e4c2",
   464 => x"f1c248bf",
   465 => x"ecc258c0",
   466 => x"c202bfd0",
   467 => x"e5c287d3",
   468 => x"e1c04ada",
   469 => x"4bc849e8",
   470 => x"7087cbe6",
   471 => x"c5c00298",
   472 => x"c348c087",
   473 => x"ecc287f6",
   474 => x"c24cbfc8",
   475 => x"c25cfcf0",
   476 => x"bf97ede4",
   477 => x"c231c849",
   478 => x"bf97ece4",
   479 => x"c249a14a",
   480 => x"bf97eee4",
   481 => x"7232d04a",
   482 => x"e4c249a1",
   483 => x"4abf97ef",
   484 => x"a17232d8",
   485 => x"c4f1c249",
   486 => x"fcf0c259",
   487 => x"f0c291bf",
   488 => x"c281bfe8",
   489 => x"c259f0f0",
   490 => x"bf97f5e4",
   491 => x"c232c84a",
   492 => x"bf97f4e4",
   493 => x"c24aa24b",
   494 => x"bf97f6e4",
   495 => x"7333d04b",
   496 => x"e4c24aa2",
   497 => x"4bbf97f7",
   498 => x"33d89bcf",
   499 => x"c24aa273",
   500 => x"c25af4f0",
   501 => x"c292748a",
   502 => x"7248f4f0",
   503 => x"c7c178a1",
   504 => x"dae4c287",
   505 => x"c849bf97",
   506 => x"d9e4c231",
   507 => x"a14abf97",
   508 => x"c731c549",
   509 => x"29c981ff",
   510 => x"59fcf0c2",
   511 => x"97dfe4c2",
   512 => x"32c84abf",
   513 => x"97dee4c2",
   514 => x"4aa24bbf",
   515 => x"5ac4f1c2",
   516 => x"bffcf0c2",
   517 => x"c2826e92",
   518 => x"c25af8f0",
   519 => x"c048f0f0",
   520 => x"ecf0c278",
   521 => x"78a17248",
   522 => x"48c4f1c2",
   523 => x"bff0f0c2",
   524 => x"c8f1c278",
   525 => x"f4f0c248",
   526 => x"ecc278bf",
   527 => x"c002bfd0",
   528 => x"487487c9",
   529 => x"7e7030c4",
   530 => x"c287c9c0",
   531 => x"48bff8f0",
   532 => x"7e7030c4",
   533 => x"48d4ecc2",
   534 => x"48c1786e",
   535 => x"4d268efc",
   536 => x"4b264c26",
   537 => x"00004f26",
   538 => x"33544146",
   539 => x"20202032",
   540 => x"00000000",
   541 => x"31544146",
   542 => x"20202036",
   543 => x"00000000",
   544 => x"33544146",
   545 => x"20202032",
   546 => x"00000000",
   547 => x"33544146",
   548 => x"20202032",
   549 => x"00000000",
   550 => x"31544146",
   551 => x"20202036",
   552 => x"5b5e0e00",
   553 => x"710e5d5c",
   554 => x"d0ecc24a",
   555 => x"87cb02bf",
   556 => x"2bc74b72",
   557 => x"ffc14d72",
   558 => x"7287c99d",
   559 => x"722bc84b",
   560 => x"9dffc34d",
   561 => x"bfe8f0c2",
   562 => x"e8f9c083",
   563 => x"d902abbf",
   564 => x"ecf9c087",
   565 => x"c8e4c25b",
   566 => x"ef49731e",
   567 => x"86c487f8",
   568 => x"c5059870",
   569 => x"c048c087",
   570 => x"ecc287e6",
   571 => x"d202bfd0",
   572 => x"c4497587",
   573 => x"c8e4c291",
   574 => x"cf4c6981",
   575 => x"ffffffff",
   576 => x"7587cb9c",
   577 => x"c291c249",
   578 => x"9f81c8e4",
   579 => x"48744c69",
   580 => x"4c264d26",
   581 => x"4f264b26",
   582 => x"5c5b5e0e",
   583 => x"86f40e5d",
   584 => x"c459a6c8",
   585 => x"80c84866",
   586 => x"c0487e70",
   587 => x"49c11e78",
   588 => x"87f9cc49",
   589 => x"4c7086c4",
   590 => x"fcc0029c",
   591 => x"d8ecc287",
   592 => x"4966dc4a",
   593 => x"87c3deff",
   594 => x"c0029870",
   595 => x"4a7487eb",
   596 => x"cb4966dc",
   597 => x"cddeff4b",
   598 => x"02987087",
   599 => x"1ec087db",
   600 => x"c4029c74",
   601 => x"c24dc087",
   602 => x"754dc187",
   603 => x"87fdcb49",
   604 => x"4c7086c4",
   605 => x"c4ff059c",
   606 => x"029c7487",
   607 => x"dc87f4c1",
   608 => x"486e49a4",
   609 => x"a4da7869",
   610 => x"4d66c449",
   611 => x"699f85c4",
   612 => x"d0ecc27d",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"6d48496e",
   620 => x"c47d7080",
   621 => x"78c04866",
   622 => x"cc4966c4",
   623 => x"c4796d81",
   624 => x"81d04966",
   625 => x"a6c879c0",
   626 => x"c878c048",
   627 => x"66c44c66",
   628 => x"7482d44a",
   629 => x"7291c849",
   630 => x"41c049a1",
   631 => x"84c1796d",
   632 => x"04acb7c6",
   633 => x"c487e7ff",
   634 => x"c4c14966",
   635 => x"c179c081",
   636 => x"c087c248",
   637 => x"268ef448",
   638 => x"264c264d",
   639 => x"0e4f264b",
   640 => x"5d5c5b5e",
   641 => x"d04c710e",
   642 => x"6c4a4d66",
   643 => x"4da17249",
   644 => x"ccecc2b9",
   645 => x"baff4abf",
   646 => x"99719972",
   647 => x"87e4c002",
   648 => x"6b4ba4c4",
   649 => x"87f9f949",
   650 => x"ecc27b70",
   651 => x"6c49bfc8",
   652 => x"757c7181",
   653 => x"ccecc2b9",
   654 => x"baff4abf",
   655 => x"99719972",
   656 => x"87dcff05",
   657 => x"4d267c75",
   658 => x"4b264c26",
   659 => x"731e4f26",
   660 => x"c24b711e",
   661 => x"49bfecf0",
   662 => x"6a4aa3c4",
   663 => x"c28ac24a",
   664 => x"92bfc8ec",
   665 => x"c249a172",
   666 => x"4abfccec",
   667 => x"a1729a6b",
   668 => x"ecf9c049",
   669 => x"1e66c859",
   670 => x"87dae971",
   671 => x"987086c4",
   672 => x"c087c405",
   673 => x"c187c248",
   674 => x"264b2648",
   675 => x"1e731e4f",
   676 => x"f0c24b71",
   677 => x"c449bfec",
   678 => x"4a6a4aa3",
   679 => x"ecc28ac2",
   680 => x"7292bfc8",
   681 => x"ecc249a1",
   682 => x"6b4abfcc",
   683 => x"49a1729a",
   684 => x"59ecf9c0",
   685 => x"711e66c8",
   686 => x"c487c6e5",
   687 => x"05987086",
   688 => x"48c087c4",
   689 => x"48c187c2",
   690 => x"4f264b26",
   691 => x"5c5b5e0e",
   692 => x"86e00e5d",
   693 => x"f0c04b71",
   694 => x"29c94966",
   695 => x"c259a6c8",
   696 => x"49bfccec",
   697 => x"4a71b9ff",
   698 => x"d89a66c4",
   699 => x"996b5aa6",
   700 => x"c459a6d0",
   701 => x"a6d07ea3",
   702 => x"78bf6e48",
   703 => x"cc4866d4",
   704 => x"c605a866",
   705 => x"7b66c487",
   706 => x"d887c1c3",
   707 => x"ffc148a6",
   708 => x"ffffffff",
   709 => x"ff80c478",
   710 => x"c84cc078",
   711 => x"a3d448a6",
   712 => x"c8497478",
   713 => x"8166c891",
   714 => x"4d4a66d4",
   715 => x"b7c08d69",
   716 => x"87ce04ad",
   717 => x"adb766d8",
   718 => x"c087c703",
   719 => x"dc5ca6e0",
   720 => x"84c15da6",
   721 => x"04acb7c6",
   722 => x"dc87d0ff",
   723 => x"b7c04866",
   724 => x"87d004a8",
   725 => x"c84966dc",
   726 => x"8166c891",
   727 => x"486e7b21",
   728 => x"87c97869",
   729 => x"a3cc7bc0",
   730 => x"69486e49",
   731 => x"4866c478",
   732 => x"a6c8886b",
   733 => x"c8ecc258",
   734 => x"90c848bf",
   735 => x"66c47e70",
   736 => x"01a86e48",
   737 => x"66c487c9",
   738 => x"03a86e48",
   739 => x"c187f3c0",
   740 => x"6a4aa3c4",
   741 => x"c891c849",
   742 => x"66cc8166",
   743 => x"c8496a79",
   744 => x"8166c891",
   745 => x"66d081c4",
   746 => x"487e6a79",
   747 => x"c705a8c5",
   748 => x"48a6c887",
   749 => x"87c778c0",
   750 => x"80c1486e",
   751 => x"c858a6cc",
   752 => x"66c47a66",
   753 => x"f849731e",
   754 => x"86c487f5",
   755 => x"1ec8e4c2",
   756 => x"f9f94973",
   757 => x"49a3d087",
   758 => x"7966f4c0",
   759 => x"268edcff",
   760 => x"264c264d",
   761 => x"0e4f264b",
   762 => x"0e5c5b5e",
   763 => x"4bc04a71",
   764 => x"c0029a72",
   765 => x"a2da87e0",
   766 => x"4b699f49",
   767 => x"bfd0ecc2",
   768 => x"d487cf02",
   769 => x"699f49a2",
   770 => x"ffc04c49",
   771 => x"34d09cff",
   772 => x"4cc087c2",
   773 => x"9b73b374",
   774 => x"4a87df02",
   775 => x"ecc28ac2",
   776 => x"9249bfc8",
   777 => x"bfecf0c2",
   778 => x"c2807248",
   779 => x"7158ccf1",
   780 => x"c230c448",
   781 => x"c058d8ec",
   782 => x"f0c287e9",
   783 => x"c24bbff0",
   784 => x"c248c8f1",
   785 => x"78bff4f0",
   786 => x"bfd0ecc2",
   787 => x"c287c902",
   788 => x"49bfc8ec",
   789 => x"87c731c4",
   790 => x"bff8f0c2",
   791 => x"c231c449",
   792 => x"c259d8ec",
   793 => x"265bc8f1",
   794 => x"264b264c",
   795 => x"5b5e0e4f",
   796 => x"f00e5d5c",
   797 => x"59a6c886",
   798 => x"ffffffcf",
   799 => x"7ec04cf8",
   800 => x"d80266c4",
   801 => x"c4e4c287",
   802 => x"c278c048",
   803 => x"c248fce3",
   804 => x"78bfc8f1",
   805 => x"48c0e4c2",
   806 => x"bfc4f1c2",
   807 => x"e5ecc278",
   808 => x"c250c048",
   809 => x"49bfd4ec",
   810 => x"bfc4e4c2",
   811 => x"03aa714a",
   812 => x"7287ccc4",
   813 => x"0599cf49",
   814 => x"c087eac0",
   815 => x"c248e8f9",
   816 => x"78bffce3",
   817 => x"1ec8e4c2",
   818 => x"bffce3c2",
   819 => x"fce3c249",
   820 => x"78a1c148",
   821 => x"fddfff71",
   822 => x"c086c487",
   823 => x"c248e4f9",
   824 => x"cc78c8e4",
   825 => x"e4f9c087",
   826 => x"e0c048bf",
   827 => x"e8f9c080",
   828 => x"c4e4c258",
   829 => x"80c148bf",
   830 => x"58c8e4c2",
   831 => x"000e6427",
   832 => x"bf97bf00",
   833 => x"c2029d4d",
   834 => x"e5c387e5",
   835 => x"dec202ad",
   836 => x"e4f9c087",
   837 => x"a3cb4bbf",
   838 => x"cf4c1149",
   839 => x"d2c105ac",
   840 => x"df497587",
   841 => x"cd89c199",
   842 => x"d8ecc291",
   843 => x"4aa3c181",
   844 => x"a3c35112",
   845 => x"c551124a",
   846 => x"51124aa3",
   847 => x"124aa3c7",
   848 => x"4aa3c951",
   849 => x"a3ce5112",
   850 => x"d051124a",
   851 => x"51124aa3",
   852 => x"124aa3d2",
   853 => x"4aa3d451",
   854 => x"a3d65112",
   855 => x"d851124a",
   856 => x"51124aa3",
   857 => x"124aa3dc",
   858 => x"4aa3de51",
   859 => x"7ec15112",
   860 => x"7487fcc0",
   861 => x"0599c849",
   862 => x"7487edc0",
   863 => x"0599d049",
   864 => x"e0c087d3",
   865 => x"ccc00266",
   866 => x"c0497387",
   867 => x"700f66e0",
   868 => x"d3c00298",
   869 => x"c0056e87",
   870 => x"ecc287c6",
   871 => x"50c048d8",
   872 => x"bfe4f9c0",
   873 => x"87ebc248",
   874 => x"48e5ecc2",
   875 => x"c27e50c0",
   876 => x"49bfd4ec",
   877 => x"bfc4e4c2",
   878 => x"04aa714a",
   879 => x"cf87f4fb",
   880 => x"f8ffffff",
   881 => x"c8f1c24c",
   882 => x"c8c005bf",
   883 => x"d0ecc287",
   884 => x"fcc102bf",
   885 => x"c0e4c287",
   886 => x"c4eb49bf",
   887 => x"c4e4c287",
   888 => x"48a6c458",
   889 => x"bfc0e4c2",
   890 => x"d0ecc278",
   891 => x"dbc002bf",
   892 => x"4966c487",
   893 => x"a9749974",
   894 => x"87c8c002",
   895 => x"c048a6c8",
   896 => x"87e7c078",
   897 => x"c148a6c8",
   898 => x"87dfc078",
   899 => x"cf4966c4",
   900 => x"a999f8ff",
   901 => x"87c8c002",
   902 => x"c048a6cc",
   903 => x"87c5c078",
   904 => x"c148a6cc",
   905 => x"48a6c878",
   906 => x"c87866cc",
   907 => x"e0c00566",
   908 => x"4966c487",
   909 => x"ecc289c2",
   910 => x"914abfc8",
   911 => x"bfecf0c2",
   912 => x"fce3c24a",
   913 => x"78a17248",
   914 => x"48c4e4c2",
   915 => x"d2f978c0",
   916 => x"cf48c087",
   917 => x"f8ffffff",
   918 => x"268ef04c",
   919 => x"264c264d",
   920 => x"004f264b",
   921 => x"00000000",
   922 => x"ffffffff",
   923 => x"48d4ff1e",
   924 => x"6878ffc3",
   925 => x"1e4f2648",
   926 => x"c348d4ff",
   927 => x"d0ff78ff",
   928 => x"78e1c048",
   929 => x"d448d4ff",
   930 => x"1e4f2678",
   931 => x"c048d0ff",
   932 => x"4f2678e0",
   933 => x"87d4ff1e",
   934 => x"02994970",
   935 => x"fbc087c6",
   936 => x"87f105a9",
   937 => x"4f264871",
   938 => x"5c5b5e0e",
   939 => x"c04b710e",
   940 => x"87f8fe4c",
   941 => x"02994970",
   942 => x"c087f9c0",
   943 => x"c002a9ec",
   944 => x"fbc087f2",
   945 => x"ebc002a9",
   946 => x"b766cc87",
   947 => x"87c703ac",
   948 => x"c20266d0",
   949 => x"71537187",
   950 => x"87c20299",
   951 => x"cbfe84c1",
   952 => x"99497087",
   953 => x"c087cd02",
   954 => x"c702a9ec",
   955 => x"a9fbc087",
   956 => x"87d5ff05",
   957 => x"c30266d0",
   958 => x"7b97c087",
   959 => x"05a9fbc0",
   960 => x"4a7487c7",
   961 => x"c28a0ac0",
   962 => x"724a7487",
   963 => x"264c2648",
   964 => x"1e4f264b",
   965 => x"7087d5fd",
   966 => x"f0c04a49",
   967 => x"87c904aa",
   968 => x"01aaf9c0",
   969 => x"f0c087c3",
   970 => x"aac1c18a",
   971 => x"c187c904",
   972 => x"c301aada",
   973 => x"8af7c087",
   974 => x"4f264872",
   975 => x"5c5b5e0e",
   976 => x"86f80e5d",
   977 => x"7ec04c71",
   978 => x"c087ecfc",
   979 => x"dcffc04b",
   980 => x"c049bf97",
   981 => x"87cf04a9",
   982 => x"c187f9fc",
   983 => x"dcffc083",
   984 => x"ab49bf97",
   985 => x"c087f106",
   986 => x"bf97dcff",
   987 => x"fb87cf02",
   988 => x"497087fa",
   989 => x"87c60299",
   990 => x"05a9ecc0",
   991 => x"4bc087f1",
   992 => x"7087e9fb",
   993 => x"87e4fb4d",
   994 => x"fb58a6c8",
   995 => x"4a7087de",
   996 => x"a4c883c1",
   997 => x"49699749",
   998 => x"87da05ad",
   999 => x"9749a4c9",
  1000 => x"66c44969",
  1001 => x"87ce05a9",
  1002 => x"9749a4ca",
  1003 => x"05aa4969",
  1004 => x"7ec187c4",
  1005 => x"ecc087d0",
  1006 => x"87c602ad",
  1007 => x"05adfbc0",
  1008 => x"4bc087c4",
  1009 => x"026e7ec1",
  1010 => x"fa87f5fe",
  1011 => x"487387fd",
  1012 => x"4d268ef8",
  1013 => x"4b264c26",
  1014 => x"00004f26",
  1015 => x"1e731e00",
  1016 => x"c84bd4ff",
  1017 => x"d0ff4a66",
  1018 => x"78c5c848",
  1019 => x"c148d4ff",
  1020 => x"7b1178d4",
  1021 => x"f9058ac1",
  1022 => x"48d0ff87",
  1023 => x"4b2678c4",
  1024 => x"5e0e4f26",
  1025 => x"0e5d5c5b",
  1026 => x"7e7186f8",
  1027 => x"f1c21e6e",
  1028 => x"c3e449dc",
  1029 => x"7086c487",
  1030 => x"e4c40298",
  1031 => x"f4ecc187",
  1032 => x"496e4cbf",
  1033 => x"c887d5fc",
  1034 => x"987058a6",
  1035 => x"c487c505",
  1036 => x"78c148a6",
  1037 => x"c548d0ff",
  1038 => x"48d4ff78",
  1039 => x"c478d5c1",
  1040 => x"89c14966",
  1041 => x"ecc131c6",
  1042 => x"4abf97ec",
  1043 => x"ffb07148",
  1044 => x"ff7808d4",
  1045 => x"78c448d0",
  1046 => x"97d8f1c2",
  1047 => x"99d049bf",
  1048 => x"c587dd02",
  1049 => x"48d4ff78",
  1050 => x"c078d6c1",
  1051 => x"48d4ff4a",
  1052 => x"c178ffc3",
  1053 => x"aae0c082",
  1054 => x"ff87f204",
  1055 => x"78c448d0",
  1056 => x"c348d4ff",
  1057 => x"d0ff78ff",
  1058 => x"ff78c548",
  1059 => x"d3c148d4",
  1060 => x"ff78c178",
  1061 => x"78c448d0",
  1062 => x"06acb7c0",
  1063 => x"c287cbc2",
  1064 => x"4bbfe4f1",
  1065 => x"737e748c",
  1066 => x"ddc1029b",
  1067 => x"4dc0c887",
  1068 => x"abb7c08b",
  1069 => x"c887c603",
  1070 => x"c04da3c0",
  1071 => x"d8f1c24b",
  1072 => x"d049bf97",
  1073 => x"87cf0299",
  1074 => x"f1c21ec0",
  1075 => x"fde549dc",
  1076 => x"7086c487",
  1077 => x"c287d84c",
  1078 => x"c21ec8e4",
  1079 => x"e549dcf1",
  1080 => x"4c7087ec",
  1081 => x"e4c21e75",
  1082 => x"f0fb49c8",
  1083 => x"7486c887",
  1084 => x"87c5059c",
  1085 => x"cac148c0",
  1086 => x"c21ec187",
  1087 => x"e349dcf1",
  1088 => x"86c487fd",
  1089 => x"fe059b73",
  1090 => x"4c6e87e3",
  1091 => x"06acb7c0",
  1092 => x"f1c287d1",
  1093 => x"78c048dc",
  1094 => x"78c080d0",
  1095 => x"f1c280f4",
  1096 => x"c078bfe8",
  1097 => x"fd01acb7",
  1098 => x"d0ff87f5",
  1099 => x"ff78c548",
  1100 => x"d3c148d4",
  1101 => x"ff78c078",
  1102 => x"78c448d0",
  1103 => x"c2c048c1",
  1104 => x"f848c087",
  1105 => x"264d268e",
  1106 => x"264b264c",
  1107 => x"5b5e0e4f",
  1108 => x"fc0e5d5c",
  1109 => x"c04d7186",
  1110 => x"04ad4c4b",
  1111 => x"c087e8c0",
  1112 => x"741efcfc",
  1113 => x"87c4029c",
  1114 => x"87c24ac0",
  1115 => x"49724ac1",
  1116 => x"c487faeb",
  1117 => x"c17e7086",
  1118 => x"c2056e83",
  1119 => x"c14b7587",
  1120 => x"06ab7584",
  1121 => x"6e87d8ff",
  1122 => x"268efc48",
  1123 => x"264c264d",
  1124 => x"0e4f264b",
  1125 => x"0e5c5b5e",
  1126 => x"66cc4b71",
  1127 => x"4c87d802",
  1128 => x"028cf0c0",
  1129 => x"4a7487d8",
  1130 => x"d1028ac1",
  1131 => x"cd028a87",
  1132 => x"c9028a87",
  1133 => x"7387d987",
  1134 => x"87c6f949",
  1135 => x"1e7487d2",
  1136 => x"d9c149c0",
  1137 => x"1e7487ca",
  1138 => x"d9c14973",
  1139 => x"86c887c2",
  1140 => x"4b264c26",
  1141 => x"5e0e4f26",
  1142 => x"0e5d5c5b",
  1143 => x"4c7186fc",
  1144 => x"c291de49",
  1145 => x"714dfcf2",
  1146 => x"026d9785",
  1147 => x"c287dcc1",
  1148 => x"49bfecf2",
  1149 => x"fd718174",
  1150 => x"7e7087d3",
  1151 => x"c0029848",
  1152 => x"f2c287f2",
  1153 => x"4a704bf0",
  1154 => x"fbfe49cb",
  1155 => x"4b7487f2",
  1156 => x"ecc193cc",
  1157 => x"83c483f8",
  1158 => x"7bd8c9c1",
  1159 => x"c2c14974",
  1160 => x"7b7587ea",
  1161 => x"97f0ecc1",
  1162 => x"c21e49bf",
  1163 => x"fd49f0f2",
  1164 => x"86c487e1",
  1165 => x"c2c14974",
  1166 => x"49c087d2",
  1167 => x"87edc3c1",
  1168 => x"48d4f1c2",
  1169 => x"c04950c0",
  1170 => x"fc87c5e1",
  1171 => x"264d268e",
  1172 => x"264b264c",
  1173 => x"0000004f",
  1174 => x"64616f4c",
  1175 => x"2e676e69",
  1176 => x"00002e2e",
  1177 => x"61422080",
  1178 => x"00006b63",
  1179 => x"64616f4c",
  1180 => x"202e2a20",
  1181 => x"00000000",
  1182 => x"0000203a",
  1183 => x"61422080",
  1184 => x"00006b63",
  1185 => x"78452080",
  1186 => x"00007469",
  1187 => x"49204453",
  1188 => x"2e74696e",
  1189 => x"0000002e",
  1190 => x"00004b4f",
  1191 => x"544f4f42",
  1192 => x"20202020",
  1193 => x"004d4f52",
  1194 => x"711e731e",
  1195 => x"f2c2494b",
  1196 => x"7181bfec",
  1197 => x"7087d6fa",
  1198 => x"c4029a4a",
  1199 => x"e6e44987",
  1200 => x"ecf2c287",
  1201 => x"7378c048",
  1202 => x"87fac149",
  1203 => x"4f264b26",
  1204 => x"711e731e",
  1205 => x"4aa3c44b",
  1206 => x"87d0c102",
  1207 => x"dc028ac1",
  1208 => x"c0028a87",
  1209 => x"058a87f2",
  1210 => x"c287d3c1",
  1211 => x"02bfecf2",
  1212 => x"4887cbc1",
  1213 => x"f2c288c1",
  1214 => x"c1c158f0",
  1215 => x"ecf2c287",
  1216 => x"89c649bf",
  1217 => x"59f0f2c2",
  1218 => x"03a9b7c0",
  1219 => x"c287efc0",
  1220 => x"c048ecf2",
  1221 => x"87e6c078",
  1222 => x"bfe8f2c2",
  1223 => x"c287df02",
  1224 => x"48bfecf2",
  1225 => x"f2c280c1",
  1226 => x"87d258f0",
  1227 => x"bfe8f2c2",
  1228 => x"c287cb02",
  1229 => x"48bfecf2",
  1230 => x"f2c280c6",
  1231 => x"497358f0",
  1232 => x"4b2687c4",
  1233 => x"5e0e4f26",
  1234 => x"0e5d5c5b",
  1235 => x"a6d086f0",
  1236 => x"c8e4c259",
  1237 => x"c24cc04d",
  1238 => x"c148e8f2",
  1239 => x"48a6c478",
  1240 => x"7e7578c0",
  1241 => x"bfecf2c2",
  1242 => x"06a8c048",
  1243 => x"7587fac0",
  1244 => x"c8e4c27e",
  1245 => x"c0029848",
  1246 => x"fcc087ef",
  1247 => x"66c81efc",
  1248 => x"c087c402",
  1249 => x"c187c24d",
  1250 => x"e349754d",
  1251 => x"86c487df",
  1252 => x"84c17e70",
  1253 => x"c14866c4",
  1254 => x"58a6c880",
  1255 => x"bfecf2c2",
  1256 => x"87c503ac",
  1257 => x"d1ff056e",
  1258 => x"c04d6e87",
  1259 => x"029d754c",
  1260 => x"c087e0c3",
  1261 => x"c81efcfc",
  1262 => x"87c70266",
  1263 => x"c048a6cc",
  1264 => x"cc87c578",
  1265 => x"78c148a6",
  1266 => x"e24966cc",
  1267 => x"86c487df",
  1268 => x"98487e70",
  1269 => x"87e8c202",
  1270 => x"9781cb49",
  1271 => x"99d04969",
  1272 => x"87d6c102",
  1273 => x"4ae8cac1",
  1274 => x"91cc4974",
  1275 => x"81f8ecc1",
  1276 => x"81c87972",
  1277 => x"7451ffc3",
  1278 => x"c291de49",
  1279 => x"714dfcf2",
  1280 => x"97c1c285",
  1281 => x"49a5c17d",
  1282 => x"c251e0c0",
  1283 => x"bf97d8ec",
  1284 => x"c187d202",
  1285 => x"4ba5c284",
  1286 => x"4ad8ecc2",
  1287 => x"f3fe49db",
  1288 => x"dbc187de",
  1289 => x"49a5cd87",
  1290 => x"84c151c0",
  1291 => x"6e4ba5c2",
  1292 => x"fe49cb4a",
  1293 => x"c187c9f3",
  1294 => x"c7c187c6",
  1295 => x"49744ad6",
  1296 => x"ecc191cc",
  1297 => x"797281f8",
  1298 => x"97d8ecc2",
  1299 => x"87d802bf",
  1300 => x"91de4974",
  1301 => x"f2c284c1",
  1302 => x"83714bfc",
  1303 => x"4ad8ecc2",
  1304 => x"f2fe49dd",
  1305 => x"87d887da",
  1306 => x"93de4b74",
  1307 => x"83fcf2c2",
  1308 => x"c049a3cb",
  1309 => x"7384c151",
  1310 => x"49cb4a6e",
  1311 => x"87c0f2fe",
  1312 => x"c14866c4",
  1313 => x"58a6c880",
  1314 => x"c003acc7",
  1315 => x"056e87c5",
  1316 => x"c787e0fc",
  1317 => x"e6c003ac",
  1318 => x"e8f2c287",
  1319 => x"c178c048",
  1320 => x"744ad6c7",
  1321 => x"c191cc49",
  1322 => x"7281f8ec",
  1323 => x"de497479",
  1324 => x"fcf2c291",
  1325 => x"c151c081",
  1326 => x"04acc784",
  1327 => x"c187daff",
  1328 => x"c048d4ee",
  1329 => x"c180f750",
  1330 => x"c140ecd4",
  1331 => x"c878e4c9",
  1332 => x"d0cbc180",
  1333 => x"4966cc78",
  1334 => x"87f0f7c0",
  1335 => x"4d268ef0",
  1336 => x"4b264c26",
  1337 => x"731e4f26",
  1338 => x"494b711e",
  1339 => x"ecc191cc",
  1340 => x"a1c881f8",
  1341 => x"ececc14a",
  1342 => x"c9501248",
  1343 => x"ffc04aa1",
  1344 => x"501248dc",
  1345 => x"ecc181ca",
  1346 => x"501148f0",
  1347 => x"97f0ecc1",
  1348 => x"c01e49bf",
  1349 => x"87fbf149",
  1350 => x"e9f84973",
  1351 => x"268efc87",
  1352 => x"1e4f264b",
  1353 => x"f8c049c0",
  1354 => x"4f2687c3",
  1355 => x"494a711e",
  1356 => x"ecc191cc",
  1357 => x"81c881f8",
  1358 => x"48d4f1c2",
  1359 => x"f0c05011",
  1360 => x"edfe49a2",
  1361 => x"49c087c6",
  1362 => x"2687c5d5",
  1363 => x"d4ff1e4f",
  1364 => x"7affc34a",
  1365 => x"c048d0ff",
  1366 => x"7ade78e1",
  1367 => x"c8487a71",
  1368 => x"7a7028b7",
  1369 => x"b7d04871",
  1370 => x"717a7028",
  1371 => x"28b7d848",
  1372 => x"d0ff7a70",
  1373 => x"78e0c048",
  1374 => x"5e0e4f26",
  1375 => x"0e5d5c5b",
  1376 => x"4d7186f4",
  1377 => x"c191cc49",
  1378 => x"c881f8ec",
  1379 => x"a1ca4aa1",
  1380 => x"48a6c47e",
  1381 => x"bfd0f1c2",
  1382 => x"bf976e78",
  1383 => x"4c66c44b",
  1384 => x"48122c73",
  1385 => x"7058a6cc",
  1386 => x"c984c19c",
  1387 => x"49699781",
  1388 => x"c204acb7",
  1389 => x"6e4cc087",
  1390 => x"c84abf97",
  1391 => x"31724966",
  1392 => x"66c4b9ff",
  1393 => x"72487499",
  1394 => x"b14a7030",
  1395 => x"59d4f1c2",
  1396 => x"87f9fd71",
  1397 => x"f2c21ec7",
  1398 => x"c11ebfe4",
  1399 => x"c21ef8ec",
  1400 => x"bf97d4f1",
  1401 => x"87f4c149",
  1402 => x"f3c04975",
  1403 => x"8ee887de",
  1404 => x"4c264d26",
  1405 => x"4f264b26",
  1406 => x"711e731e",
  1407 => x"f9fd494b",
  1408 => x"fd497387",
  1409 => x"4b2687f4",
  1410 => x"731e4f26",
  1411 => x"c24b711e",
  1412 => x"d6024aa3",
  1413 => x"058ac187",
  1414 => x"c287e2c0",
  1415 => x"02bfe4f2",
  1416 => x"c14887db",
  1417 => x"e8f2c288",
  1418 => x"c287d258",
  1419 => x"02bfe8f2",
  1420 => x"f2c287cb",
  1421 => x"c148bfe4",
  1422 => x"e8f2c280",
  1423 => x"c21ec758",
  1424 => x"1ebfe4f2",
  1425 => x"1ef8ecc1",
  1426 => x"97d4f1c2",
  1427 => x"87cc49bf",
  1428 => x"f1c04973",
  1429 => x"8ef487f6",
  1430 => x"4f264b26",
  1431 => x"5c5b5e0e",
  1432 => x"ccff0e5d",
  1433 => x"a6e8c086",
  1434 => x"48a6cc59",
  1435 => x"80c478c0",
  1436 => x"80c478c0",
  1437 => x"80c478c0",
  1438 => x"7866c8c1",
  1439 => x"78c180c4",
  1440 => x"78c180c4",
  1441 => x"48e8f2c2",
  1442 => x"dfff78c1",
  1443 => x"c3e087e9",
  1444 => x"d7dfff87",
  1445 => x"c04d7087",
  1446 => x"c102adfb",
  1447 => x"e4c087f3",
  1448 => x"e8c10566",
  1449 => x"66c4c187",
  1450 => x"6a82c44a",
  1451 => x"ecc9c17e",
  1452 => x"20496e48",
  1453 => x"10412041",
  1454 => x"66c4c151",
  1455 => x"e6d3c148",
  1456 => x"c7496a78",
  1457 => x"c1517581",
  1458 => x"c84966c4",
  1459 => x"dc51c181",
  1460 => x"78c248a6",
  1461 => x"4966c4c1",
  1462 => x"51c081c9",
  1463 => x"4966c4c1",
  1464 => x"51c081ca",
  1465 => x"1ed81ec1",
  1466 => x"81c8496a",
  1467 => x"87f8deff",
  1468 => x"c8c186c8",
  1469 => x"a8c04866",
  1470 => x"d487c701",
  1471 => x"78c148a6",
  1472 => x"c8c187cf",
  1473 => x"88c14866",
  1474 => x"c458a6dc",
  1475 => x"c3deff87",
  1476 => x"029d7587",
  1477 => x"d487f1cb",
  1478 => x"ccc14866",
  1479 => x"cb03a866",
  1480 => x"7ec087e6",
  1481 => x"87c4ddff",
  1482 => x"c1484d70",
  1483 => x"a6c888c6",
  1484 => x"02987058",
  1485 => x"4887d6c1",
  1486 => x"a6c888c9",
  1487 => x"02987058",
  1488 => x"4887d7c5",
  1489 => x"a6c888c1",
  1490 => x"02987058",
  1491 => x"4887f8c2",
  1492 => x"a6c888c3",
  1493 => x"02987058",
  1494 => x"c14887cf",
  1495 => x"58a6c888",
  1496 => x"c4029870",
  1497 => x"fec987f4",
  1498 => x"7ef0c087",
  1499 => x"87fcdbff",
  1500 => x"ecc04d70",
  1501 => x"87c202ad",
  1502 => x"ecc07e75",
  1503 => x"87cd02ad",
  1504 => x"87e8dbff",
  1505 => x"ecc04d70",
  1506 => x"f3ff05ad",
  1507 => x"66e4c087",
  1508 => x"87eac105",
  1509 => x"02adecc0",
  1510 => x"dbff87c4",
  1511 => x"1ec087ce",
  1512 => x"66dc1eca",
  1513 => x"c193cc4b",
  1514 => x"c48366cc",
  1515 => x"496c4ca3",
  1516 => x"87f4dbff",
  1517 => x"1ede1ec1",
  1518 => x"dbff496c",
  1519 => x"86d087ea",
  1520 => x"7be6d3c1",
  1521 => x"dc49a3c8",
  1522 => x"a3c95166",
  1523 => x"66e0c049",
  1524 => x"49a3ca51",
  1525 => x"66dc516e",
  1526 => x"c080c148",
  1527 => x"d458a6e0",
  1528 => x"66d84866",
  1529 => x"87cb04a8",
  1530 => x"c14866d4",
  1531 => x"58a6d880",
  1532 => x"d887fac7",
  1533 => x"88c14866",
  1534 => x"c758a6dc",
  1535 => x"daff87ef",
  1536 => x"4d7087d2",
  1537 => x"ff87e6c7",
  1538 => x"d087c8dc",
  1539 => x"66d058a6",
  1540 => x"87c606a8",
  1541 => x"cc48a6d0",
  1542 => x"dbff7866",
  1543 => x"ecc087f5",
  1544 => x"f5c105a8",
  1545 => x"66e4c087",
  1546 => x"87e5c105",
  1547 => x"cc4966d4",
  1548 => x"66c4c191",
  1549 => x"4aa1c481",
  1550 => x"a1c84c6a",
  1551 => x"5266cc4a",
  1552 => x"79ecd4c1",
  1553 => x"87e4d8ff",
  1554 => x"029d4d70",
  1555 => x"fbc087da",
  1556 => x"87d402ad",
  1557 => x"d8ff5475",
  1558 => x"4d7087d2",
  1559 => x"c7c0029d",
  1560 => x"adfbc087",
  1561 => x"87ecff05",
  1562 => x"c254e0c0",
  1563 => x"97c054c1",
  1564 => x"4866d47c",
  1565 => x"04a866d8",
  1566 => x"d487cbc0",
  1567 => x"80c14866",
  1568 => x"c558a6d8",
  1569 => x"66d887e7",
  1570 => x"dc88c148",
  1571 => x"dcc558a6",
  1572 => x"ffd7ff87",
  1573 => x"c54d7087",
  1574 => x"66cc87d3",
  1575 => x"66e4c048",
  1576 => x"f4c405a8",
  1577 => x"a6e8c087",
  1578 => x"ff78c048",
  1579 => x"7087e4d9",
  1580 => x"ded9ff7e",
  1581 => x"a6f0c087",
  1582 => x"a8ecc058",
  1583 => x"87c7c005",
  1584 => x"786e48a6",
  1585 => x"ff87c4c0",
  1586 => x"d487e1d6",
  1587 => x"91cc4966",
  1588 => x"4866c4c1",
  1589 => x"a6c88071",
  1590 => x"4a66c458",
  1591 => x"66c482c8",
  1592 => x"6e81ca49",
  1593 => x"66ecc051",
  1594 => x"6e81c149",
  1595 => x"7148c189",
  1596 => x"c1497030",
  1597 => x"7a977189",
  1598 => x"bfd0f1c2",
  1599 => x"97296e49",
  1600 => x"71484a6a",
  1601 => x"a6f4c098",
  1602 => x"4866c458",
  1603 => x"a6cc80c4",
  1604 => x"bf66c858",
  1605 => x"66e4c04c",
  1606 => x"a866cc48",
  1607 => x"87c5c002",
  1608 => x"c2c07ec0",
  1609 => x"6e7ec187",
  1610 => x"1ee0c01e",
  1611 => x"d5ff4974",
  1612 => x"86c887f6",
  1613 => x"b7c04d70",
  1614 => x"d4c106ad",
  1615 => x"c8847587",
  1616 => x"c049bf66",
  1617 => x"897481e0",
  1618 => x"f8c9c14b",
  1619 => x"defe714a",
  1620 => x"84c287ee",
  1621 => x"e8c07e74",
  1622 => x"80c14866",
  1623 => x"58a6ecc0",
  1624 => x"4966f0c0",
  1625 => x"a97081c1",
  1626 => x"87c5c002",
  1627 => x"c2c04cc0",
  1628 => x"744cc187",
  1629 => x"bf66cc1e",
  1630 => x"81e0c049",
  1631 => x"718966c4",
  1632 => x"4966c81e",
  1633 => x"87e0d4ff",
  1634 => x"b7c086c8",
  1635 => x"c5ff01a8",
  1636 => x"66e8c087",
  1637 => x"87d3c002",
  1638 => x"c94966c4",
  1639 => x"66e8c081",
  1640 => x"4866c451",
  1641 => x"78fad5c1",
  1642 => x"c487cec0",
  1643 => x"81c94966",
  1644 => x"66c451c2",
  1645 => x"f8d7c148",
  1646 => x"4866d478",
  1647 => x"04a866d8",
  1648 => x"d487cbc0",
  1649 => x"80c14866",
  1650 => x"c058a6d8",
  1651 => x"66d887d1",
  1652 => x"dc88c148",
  1653 => x"c6c058a6",
  1654 => x"f7d2ff87",
  1655 => x"cc4d7087",
  1656 => x"78c048a6",
  1657 => x"ff87c6c0",
  1658 => x"7087e9d2",
  1659 => x"66e0c04d",
  1660 => x"c080c148",
  1661 => x"7558a6e4",
  1662 => x"cbc0029d",
  1663 => x"4866d487",
  1664 => x"a866ccc1",
  1665 => x"87daf404",
  1666 => x"c74866d4",
  1667 => x"e1c003a8",
  1668 => x"4c66d487",
  1669 => x"48e8f2c2",
  1670 => x"497478c0",
  1671 => x"c4c191cc",
  1672 => x"a1c48166",
  1673 => x"c04a6a4a",
  1674 => x"84c17952",
  1675 => x"ff04acc7",
  1676 => x"e4c087e2",
  1677 => x"e2c00266",
  1678 => x"66c4c187",
  1679 => x"81d4c149",
  1680 => x"4a66c4c1",
  1681 => x"c082dcc1",
  1682 => x"ecd4c152",
  1683 => x"66c4c179",
  1684 => x"81d8c149",
  1685 => x"79fcc9c1",
  1686 => x"c187d6c0",
  1687 => x"c14966c4",
  1688 => x"c4c181d4",
  1689 => x"d8c14a66",
  1690 => x"c4cac182",
  1691 => x"e3d4c17a",
  1692 => x"cad8c179",
  1693 => x"66c4c14a",
  1694 => x"81e0c149",
  1695 => x"d0ff7972",
  1696 => x"66d087c9",
  1697 => x"8eccff48",
  1698 => x"4c264d26",
  1699 => x"4f264b26",
  1700 => x"c21ec71e",
  1701 => x"1ebfe4f2",
  1702 => x"1ef8ecc1",
  1703 => x"97d4f1c2",
  1704 => x"f7ee49bf",
  1705 => x"f8ecc187",
  1706 => x"ede1c049",
  1707 => x"268ef487",
  1708 => x"1e731e4f",
  1709 => x"c287cfc7",
  1710 => x"c048f0f2",
  1711 => x"48d4ff50",
  1712 => x"c178ffc3",
  1713 => x"fe49ccca",
  1714 => x"fe87dcd7",
  1715 => x"7087f1e2",
  1716 => x"87cd0298",
  1717 => x"87cfecfe",
  1718 => x"c4029870",
  1719 => x"c24ac187",
  1720 => x"724ac087",
  1721 => x"87c8029a",
  1722 => x"49d8cac1",
  1723 => x"87f7d6fe",
  1724 => x"48e4f2c2",
  1725 => x"f1c278c0",
  1726 => x"50c048d4",
  1727 => x"87d0fe49",
  1728 => x"87f1f6c0",
  1729 => x"029b4b70",
  1730 => x"eec187cf",
  1731 => x"49c75bd4",
  1732 => x"c187f9de",
  1733 => x"d4e0c049",
  1734 => x"87f3c287",
  1735 => x"87dae1c0",
  1736 => x"87f5efc0",
  1737 => x"2687f5ff",
  1738 => x"004f264b",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"00000001",
  1742 => x"000011d6",
  1743 => x"00002cbc",
  1744 => x"00000000",
  1745 => x"000011d6",
  1746 => x"00002cda",
  1747 => x"00000000",
  1748 => x"000011d6",
  1749 => x"00002cf8",
  1750 => x"00000000",
  1751 => x"000011d6",
  1752 => x"00002d16",
  1753 => x"00000000",
  1754 => x"000011d6",
  1755 => x"00002d34",
  1756 => x"00000000",
  1757 => x"000011d6",
  1758 => x"00002d52",
  1759 => x"00000000",
  1760 => x"000011d6",
  1761 => x"00002d70",
  1762 => x"00000000",
  1763 => x"0000152c",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"000012d0",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"0000129c",
  1770 => x"db86fc1e",
  1771 => x"fc7e7087",
  1772 => x"1e4f268e",
  1773 => x"c048f0fe",
  1774 => x"7909cd78",
  1775 => x"1e4f2609",
  1776 => x"49e8eec1",
  1777 => x"4f2687ed",
  1778 => x"bff0fe1e",
  1779 => x"1e4f2648",
  1780 => x"c148f0fe",
  1781 => x"1e4f2678",
  1782 => x"c048f0fe",
  1783 => x"1e4f2678",
  1784 => x"52c04a71",
  1785 => x"0e4f2651",
  1786 => x"5d5c5b5e",
  1787 => x"7186f40e",
  1788 => x"7e6d974d",
  1789 => x"974ca5c1",
  1790 => x"a6c8486c",
  1791 => x"c4486e58",
  1792 => x"c505a866",
  1793 => x"c048ff87",
  1794 => x"caff87e6",
  1795 => x"49a5c287",
  1796 => x"714b6c97",
  1797 => x"6b974ba3",
  1798 => x"7e6c974b",
  1799 => x"80c1486e",
  1800 => x"c758a6c8",
  1801 => x"58a6cc98",
  1802 => x"fe7c9770",
  1803 => x"487387e1",
  1804 => x"4d268ef4",
  1805 => x"4b264c26",
  1806 => x"731e4f26",
  1807 => x"fe86f41e",
  1808 => x"bfe087d5",
  1809 => x"e0c0494b",
  1810 => x"c00299c0",
  1811 => x"4a7387ea",
  1812 => x"c29affc3",
  1813 => x"bf97e4f6",
  1814 => x"e6f6c249",
  1815 => x"c2517281",
  1816 => x"bf97e4f6",
  1817 => x"c1486e7e",
  1818 => x"58a6c880",
  1819 => x"a6cc98c7",
  1820 => x"e4f6c258",
  1821 => x"5066c848",
  1822 => x"7087cdfd",
  1823 => x"87cffd7e",
  1824 => x"4b268ef4",
  1825 => x"c21e4f26",
  1826 => x"fd49e4f6",
  1827 => x"f0c187d1",
  1828 => x"defc49fa",
  1829 => x"87e8c487",
  1830 => x"5e0e4f26",
  1831 => x"0e5d5c5b",
  1832 => x"7e7186fc",
  1833 => x"c24dd4ff",
  1834 => x"fc49e4f6",
  1835 => x"4b7087f9",
  1836 => x"04abb7c0",
  1837 => x"c387f5c2",
  1838 => x"c905abf0",
  1839 => x"f8f5c187",
  1840 => x"c278c148",
  1841 => x"e0c387d6",
  1842 => x"87c905ab",
  1843 => x"48fcf5c1",
  1844 => x"c7c278c1",
  1845 => x"fcf5c187",
  1846 => x"87c602bf",
  1847 => x"4ca3c0c2",
  1848 => x"4c7387c2",
  1849 => x"bff8f5c1",
  1850 => x"87e0c002",
  1851 => x"b7c44974",
  1852 => x"f6c19129",
  1853 => x"4a7481c0",
  1854 => x"92c29acf",
  1855 => x"307248c1",
  1856 => x"baff4a70",
  1857 => x"98694872",
  1858 => x"87db7970",
  1859 => x"b7c44974",
  1860 => x"f6c19129",
  1861 => x"4a7481c0",
  1862 => x"92c29acf",
  1863 => x"307248c3",
  1864 => x"69484a70",
  1865 => x"6e7970b0",
  1866 => x"87e4c005",
  1867 => x"c848d0ff",
  1868 => x"7dc578e1",
  1869 => x"bffcf5c1",
  1870 => x"c387c302",
  1871 => x"f5c17de0",
  1872 => x"c302bff8",
  1873 => x"7df0c387",
  1874 => x"d0ff7d73",
  1875 => x"78e0c048",
  1876 => x"48fcf5c1",
  1877 => x"f5c178c0",
  1878 => x"78c048f8",
  1879 => x"49e4f6c2",
  1880 => x"7087c4fa",
  1881 => x"abb7c04b",
  1882 => x"87cbfd03",
  1883 => x"8efc48c0",
  1884 => x"4c264d26",
  1885 => x"4f264b26",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"724ac01e",
  1905 => x"c191c449",
  1906 => x"c081c0f6",
  1907 => x"d082c179",
  1908 => x"ee04aab7",
  1909 => x"0e4f2687",
  1910 => x"5d5c5b5e",
  1911 => x"f74d710e",
  1912 => x"4a7587f5",
  1913 => x"922ab7c4",
  1914 => x"82c0f6c1",
  1915 => x"9ccf4c75",
  1916 => x"496a94c2",
  1917 => x"c32b744b",
  1918 => x"7448c29b",
  1919 => x"ff4c7030",
  1920 => x"714874bc",
  1921 => x"f77a7098",
  1922 => x"487387c5",
  1923 => x"4c264d26",
  1924 => x"4f264b26",
  1925 => x"48d0ff1e",
  1926 => x"7178e1c8",
  1927 => x"08d4ff48",
  1928 => x"1e4f2678",
  1929 => x"c848d0ff",
  1930 => x"487178e1",
  1931 => x"7808d4ff",
  1932 => x"ff4866c4",
  1933 => x"267808d4",
  1934 => x"4a711e4f",
  1935 => x"1e4966c4",
  1936 => x"deff4972",
  1937 => x"48d0ff87",
  1938 => x"fc78e0c0",
  1939 => x"1e4f268e",
  1940 => x"4a711e73",
  1941 => x"abb7c24b",
  1942 => x"a387c803",
  1943 => x"ffc34a49",
  1944 => x"ce87c79a",
  1945 => x"c34a49a3",
  1946 => x"66c89aff",
  1947 => x"49721e49",
  1948 => x"fc87c6ff",
  1949 => x"264b268e",
  1950 => x"d0ff1e4f",
  1951 => x"78c9c848",
  1952 => x"d4ff4871",
  1953 => x"4f267808",
  1954 => x"494a711e",
  1955 => x"d0ff87eb",
  1956 => x"2678c848",
  1957 => x"1e731e4f",
  1958 => x"f6c24b71",
  1959 => x"c302bffc",
  1960 => x"87ebc287",
  1961 => x"c848d0ff",
  1962 => x"487378c9",
  1963 => x"ffb0e0c0",
  1964 => x"c27808d4",
  1965 => x"c048f0f6",
  1966 => x"0266c878",
  1967 => x"ffc387c5",
  1968 => x"c087c249",
  1969 => x"f8f6c249",
  1970 => x"0266cc59",
  1971 => x"d5c587c6",
  1972 => x"87c44ad5",
  1973 => x"4affffcf",
  1974 => x"5afcf6c2",
  1975 => x"48fcf6c2",
  1976 => x"4b2678c1",
  1977 => x"5e0e4f26",
  1978 => x"0e5d5c5b",
  1979 => x"f6c24d71",
  1980 => x"754bbff8",
  1981 => x"87cb029d",
  1982 => x"c191c849",
  1983 => x"714accfa",
  1984 => x"c187c482",
  1985 => x"c04accfe",
  1986 => x"7349124c",
  1987 => x"f4f6c299",
  1988 => x"b87148bf",
  1989 => x"7808d4ff",
  1990 => x"842bb7c1",
  1991 => x"04acb7c8",
  1992 => x"f6c287e7",
  1993 => x"c848bff0",
  1994 => x"f4f6c280",
  1995 => x"264d2658",
  1996 => x"264b264c",
  1997 => x"1e731e4f",
  1998 => x"4a134b71",
  1999 => x"87cb029a",
  2000 => x"e1fe4972",
  2001 => x"9a4a1387",
  2002 => x"2687f505",
  2003 => x"1e4f264b",
  2004 => x"bff0f6c2",
  2005 => x"f0f6c249",
  2006 => x"78a1c148",
  2007 => x"a9b7c0c4",
  2008 => x"ff87db03",
  2009 => x"f6c248d4",
  2010 => x"c278bff4",
  2011 => x"49bff0f6",
  2012 => x"48f0f6c2",
  2013 => x"c478a1c1",
  2014 => x"04a9b7c0",
  2015 => x"d0ff87e5",
  2016 => x"c278c848",
  2017 => x"c048fcf6",
  2018 => x"004f2678",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"5f000000",
  2022 => x"0000005f",
  2023 => x"00030300",
  2024 => x"00000303",
  2025 => x"147f7f14",
  2026 => x"00147f7f",
  2027 => x"6b2e2400",
  2028 => x"00123a6b",
  2029 => x"18366a4c",
  2030 => x"0032566c",
  2031 => x"594f7e30",
  2032 => x"40683a77",
  2033 => x"07040000",
  2034 => x"00000003",
  2035 => x"3e1c0000",
  2036 => x"00004163",
  2037 => x"63410000",
  2038 => x"00001c3e",
  2039 => x"1c3e2a08",
  2040 => x"082a3e1c",
  2041 => x"3e080800",
  2042 => x"0008083e",
  2043 => x"e0800000",
  2044 => x"00000060",
  2045 => x"08080800",
  2046 => x"00080808",
  2047 => x"60000000",
  2048 => x"00000060",
  2049 => x"18306040",
  2050 => x"0103060c",
  2051 => x"597f3e00",
  2052 => x"003e7f4d",
  2053 => x"7f060400",
  2054 => x"0000007f",
  2055 => x"71634200",
  2056 => x"00464f59",
  2057 => x"49632200",
  2058 => x"00367f49",
  2059 => x"13161c18",
  2060 => x"00107f7f",
  2061 => x"45672700",
  2062 => x"00397d45",
  2063 => x"4b7e3c00",
  2064 => x"00307949",
  2065 => x"71010100",
  2066 => x"00070f79",
  2067 => x"497f3600",
  2068 => x"00367f49",
  2069 => x"494f0600",
  2070 => x"001e3f69",
  2071 => x"66000000",
  2072 => x"00000066",
  2073 => x"e6800000",
  2074 => x"00000066",
  2075 => x"14080800",
  2076 => x"00222214",
  2077 => x"14141400",
  2078 => x"00141414",
  2079 => x"14222200",
  2080 => x"00080814",
  2081 => x"51030200",
  2082 => x"00060f59",
  2083 => x"5d417f3e",
  2084 => x"001e1f55",
  2085 => x"097f7e00",
  2086 => x"007e7f09",
  2087 => x"497f7f00",
  2088 => x"00367f49",
  2089 => x"633e1c00",
  2090 => x"00414141",
  2091 => x"417f7f00",
  2092 => x"001c3e63",
  2093 => x"497f7f00",
  2094 => x"00414149",
  2095 => x"097f7f00",
  2096 => x"00010109",
  2097 => x"417f3e00",
  2098 => x"007a7b49",
  2099 => x"087f7f00",
  2100 => x"007f7f08",
  2101 => x"7f410000",
  2102 => x"0000417f",
  2103 => x"40602000",
  2104 => x"003f7f40",
  2105 => x"1c087f7f",
  2106 => x"00416336",
  2107 => x"407f7f00",
  2108 => x"00404040",
  2109 => x"0c067f7f",
  2110 => x"007f7f06",
  2111 => x"0c067f7f",
  2112 => x"007f7f18",
  2113 => x"417f3e00",
  2114 => x"003e7f41",
  2115 => x"097f7f00",
  2116 => x"00060f09",
  2117 => x"61417f3e",
  2118 => x"00407e7f",
  2119 => x"097f7f00",
  2120 => x"00667f19",
  2121 => x"4d6f2600",
  2122 => x"00327b59",
  2123 => x"7f010100",
  2124 => x"0001017f",
  2125 => x"407f3f00",
  2126 => x"003f7f40",
  2127 => x"703f0f00",
  2128 => x"000f3f70",
  2129 => x"18307f7f",
  2130 => x"007f7f30",
  2131 => x"1c366341",
  2132 => x"4163361c",
  2133 => x"7c060301",
  2134 => x"0103067c",
  2135 => x"4d597161",
  2136 => x"00414347",
  2137 => x"7f7f0000",
  2138 => x"00004141",
  2139 => x"0c060301",
  2140 => x"40603018",
  2141 => x"41410000",
  2142 => x"00007f7f",
  2143 => x"03060c08",
  2144 => x"00080c06",
  2145 => x"80808080",
  2146 => x"00808080",
  2147 => x"03000000",
  2148 => x"00000407",
  2149 => x"54742000",
  2150 => x"00787c54",
  2151 => x"447f7f00",
  2152 => x"00387c44",
  2153 => x"447c3800",
  2154 => x"00004444",
  2155 => x"447c3800",
  2156 => x"007f7f44",
  2157 => x"547c3800",
  2158 => x"00185c54",
  2159 => x"7f7e0400",
  2160 => x"00000505",
  2161 => x"a4bc1800",
  2162 => x"007cfca4",
  2163 => x"047f7f00",
  2164 => x"00787c04",
  2165 => x"3d000000",
  2166 => x"0000407d",
  2167 => x"80808000",
  2168 => x"00007dfd",
  2169 => x"107f7f00",
  2170 => x"00446c38",
  2171 => x"3f000000",
  2172 => x"0000407f",
  2173 => x"180c7c7c",
  2174 => x"00787c0c",
  2175 => x"047c7c00",
  2176 => x"00787c04",
  2177 => x"447c3800",
  2178 => x"00387c44",
  2179 => x"24fcfc00",
  2180 => x"00183c24",
  2181 => x"243c1800",
  2182 => x"00fcfc24",
  2183 => x"047c7c00",
  2184 => x"00080c04",
  2185 => x"545c4800",
  2186 => x"00207454",
  2187 => x"7f3f0400",
  2188 => x"00004444",
  2189 => x"407c3c00",
  2190 => x"007c7c40",
  2191 => x"603c1c00",
  2192 => x"001c3c60",
  2193 => x"30607c3c",
  2194 => x"003c7c60",
  2195 => x"10386c44",
  2196 => x"00446c38",
  2197 => x"e0bc1c00",
  2198 => x"001c3c60",
  2199 => x"74644400",
  2200 => x"00444c5c",
  2201 => x"3e080800",
  2202 => x"00414177",
  2203 => x"7f000000",
  2204 => x"0000007f",
  2205 => x"77414100",
  2206 => x"0008083e",
  2207 => x"03010102",
  2208 => x"00010202",
  2209 => x"7f7f7f7f",
  2210 => x"007f7f7f",
  2211 => x"1c1c0808",
  2212 => x"7f7f3e3e",
  2213 => x"3e3e7f7f",
  2214 => x"08081c1c",
  2215 => x"7c181000",
  2216 => x"0010187c",
  2217 => x"7c301000",
  2218 => x"0010307c",
  2219 => x"60603010",
  2220 => x"00061e78",
  2221 => x"183c6642",
  2222 => x"0042663c",
  2223 => x"c26a3878",
  2224 => x"00386cc6",
  2225 => x"60000060",
  2226 => x"00600000",
  2227 => x"5c5b5e0e",
  2228 => x"86fc0e5d",
  2229 => x"f7c27e71",
  2230 => x"c04cbfc4",
  2231 => x"c41ec04b",
  2232 => x"c402ab66",
  2233 => x"c24dc087",
  2234 => x"754dc187",
  2235 => x"ee49731e",
  2236 => x"86c887e3",
  2237 => x"ef49e0c0",
  2238 => x"a4c487ec",
  2239 => x"f0496a4a",
  2240 => x"caf187f3",
  2241 => x"c184cc87",
  2242 => x"abb7c883",
  2243 => x"87cdff04",
  2244 => x"4d268efc",
  2245 => x"4b264c26",
  2246 => x"711e4f26",
  2247 => x"c8f7c24a",
  2248 => x"c8f7c25a",
  2249 => x"4978c748",
  2250 => x"2687e1fe",
  2251 => x"1e731e4f",
  2252 => x"0bfc4b71",
  2253 => x"4a730b7b",
  2254 => x"c0c19ac1",
  2255 => x"c7ed49a2",
  2256 => x"c0dac287",
  2257 => x"264b265b",
  2258 => x"4a711e4f",
  2259 => x"721e66c4",
  2260 => x"87fbeb49",
  2261 => x"4f268efc",
  2262 => x"48d4ff1e",
  2263 => x"ff78ffc3",
  2264 => x"e1c048d0",
  2265 => x"48d4ff78",
  2266 => x"487178c1",
  2267 => x"d4ff30c4",
  2268 => x"d0ff7808",
  2269 => x"78e0c048",
  2270 => x"5e0e4f26",
  2271 => x"0e5d5c5b",
  2272 => x"7ec086f4",
  2273 => x"ec48a6c8",
  2274 => x"80fc78bf",
  2275 => x"bfc4f7c2",
  2276 => x"ccf7c278",
  2277 => x"bfe84cbf",
  2278 => x"fcd9c24d",
  2279 => x"f9e349bf",
  2280 => x"e849c787",
  2281 => x"497087f1",
  2282 => x"d00599c2",
  2283 => x"f4d9c287",
  2284 => x"b9ff49bf",
  2285 => x"c19966c8",
  2286 => x"f9c10299",
  2287 => x"49e8cf87",
  2288 => x"7087fdca",
  2289 => x"e849c74b",
  2290 => x"987087cd",
  2291 => x"c887c905",
  2292 => x"99c14966",
  2293 => x"87fec002",
  2294 => x"ec48a6c8",
  2295 => x"f9e278bf",
  2296 => x"ca497387",
  2297 => x"987087e6",
  2298 => x"c287d702",
  2299 => x"49bff0d9",
  2300 => x"d9c2b9c1",
  2301 => x"fd7159f4",
  2302 => x"e8cf87de",
  2303 => x"87c0ca49",
  2304 => x"49c74b70",
  2305 => x"7087d0e7",
  2306 => x"cbff0598",
  2307 => x"4966c887",
  2308 => x"ff0599c1",
  2309 => x"d9c287c2",
  2310 => x"c14abffc",
  2311 => x"c0dac2ba",
  2312 => x"7a0afc5a",
  2313 => x"c19ac10a",
  2314 => x"e949a2c0",
  2315 => x"dac187da",
  2316 => x"87e3e649",
  2317 => x"d9c27ec1",
  2318 => x"66c848f4",
  2319 => x"fcd9c278",
  2320 => x"e9c005bf",
  2321 => x"c3497587",
  2322 => x"1e7199ff",
  2323 => x"f8fb49c0",
  2324 => x"c8497587",
  2325 => x"1e7129b7",
  2326 => x"ecfb49c1",
  2327 => x"c386c887",
  2328 => x"f2e549fd",
  2329 => x"49fac387",
  2330 => x"c787ece5",
  2331 => x"497587f4",
  2332 => x"c899ffc3",
  2333 => x"b5712db7",
  2334 => x"c0029d75",
  2335 => x"a6c887e4",
  2336 => x"bfc8ff48",
  2337 => x"4966c878",
  2338 => x"bff8d9c2",
  2339 => x"a9e0c289",
  2340 => x"87c4c003",
  2341 => x"87d04dc0",
  2342 => x"48f8d9c2",
  2343 => x"c07866c8",
  2344 => x"d9c287c6",
  2345 => x"78c048f8",
  2346 => x"99c84975",
  2347 => x"87cec005",
  2348 => x"e449f5c3",
  2349 => x"497087e1",
  2350 => x"c00299c2",
  2351 => x"f7c287e7",
  2352 => x"c002bfc8",
  2353 => x"c14887ca",
  2354 => x"ccf7c288",
  2355 => x"87d3c058",
  2356 => x"c14866c4",
  2357 => x"7e7080e0",
  2358 => x"c002bf6e",
  2359 => x"ff4b87c5",
  2360 => x"c10f7349",
  2361 => x"c449757e",
  2362 => x"cec00599",
  2363 => x"49f2c387",
  2364 => x"7087e4e3",
  2365 => x"0299c249",
  2366 => x"c287eac0",
  2367 => x"7ebfc8f7",
  2368 => x"a8b7c748",
  2369 => x"87cbc003",
  2370 => x"80c1486e",
  2371 => x"58ccf7c2",
  2372 => x"c487d0c0",
  2373 => x"e0c14a66",
  2374 => x"c0026a82",
  2375 => x"fe4b87c5",
  2376 => x"c10f7349",
  2377 => x"49fdc37e",
  2378 => x"7087ece2",
  2379 => x"0299c249",
  2380 => x"c287e6c0",
  2381 => x"02bfc8f7",
  2382 => x"c287c9c0",
  2383 => x"c048c8f7",
  2384 => x"87d3c078",
  2385 => x"c14866c4",
  2386 => x"7e7080e0",
  2387 => x"c002bf6e",
  2388 => x"fd4b87c5",
  2389 => x"c10f7349",
  2390 => x"49fac37e",
  2391 => x"7087f8e1",
  2392 => x"0299c249",
  2393 => x"c287eac0",
  2394 => x"48bfc8f7",
  2395 => x"03a8b7c7",
  2396 => x"c287c9c0",
  2397 => x"c748c8f7",
  2398 => x"87d3c078",
  2399 => x"c14866c4",
  2400 => x"7e7080e0",
  2401 => x"c002bf6e",
  2402 => x"fc4b87c5",
  2403 => x"c10f7349",
  2404 => x"c348757e",
  2405 => x"a6cc98f0",
  2406 => x"05987058",
  2407 => x"c187cec0",
  2408 => x"f2e049da",
  2409 => x"c2497087",
  2410 => x"f9c10299",
  2411 => x"49e8cf87",
  2412 => x"7087cdc3",
  2413 => x"c0f7c24b",
  2414 => x"c250c048",
  2415 => x"bf97c0f7",
  2416 => x"87d2c105",
  2417 => x"c00566c8",
  2418 => x"dac187cc",
  2419 => x"87c7e049",
  2420 => x"c1029870",
  2421 => x"bfe887c0",
  2422 => x"ffc3494d",
  2423 => x"2db7c899",
  2424 => x"daffb571",
  2425 => x"497387f4",
  2426 => x"7087e1c2",
  2427 => x"c6c00298",
  2428 => x"c0f7c287",
  2429 => x"c250c148",
  2430 => x"bf97c0f7",
  2431 => x"87d6c005",
  2432 => x"f0c34975",
  2433 => x"cdff0599",
  2434 => x"49dac187",
  2435 => x"87c7dfff",
  2436 => x"ff059870",
  2437 => x"f7c287c0",
  2438 => x"4b49bfc8",
  2439 => x"66c493cc",
  2440 => x"714b6b83",
  2441 => x"9c740f73",
  2442 => x"87e9c002",
  2443 => x"e4c0026c",
  2444 => x"ff496c87",
  2445 => x"7087e0de",
  2446 => x"0299c149",
  2447 => x"c487cbc0",
  2448 => x"f7c24ba4",
  2449 => x"6b49bfc8",
  2450 => x"84c80f4b",
  2451 => x"87c5c002",
  2452 => x"dcff056c",
  2453 => x"c0026e87",
  2454 => x"f7c287c8",
  2455 => x"f149bfc8",
  2456 => x"8ef487ea",
  2457 => x"4c264d26",
  2458 => x"4f264b26",
  2459 => x"00000010",
  2460 => x"00000000",
  2461 => x"00000000",
  2462 => x"00000000",
  2463 => x"00000000",
  2464 => x"ff4a711e",
  2465 => x"7249bfc8",
  2466 => x"4f2648a1",
  2467 => x"bfc8ff1e",
  2468 => x"c0c0fe89",
  2469 => x"a9c0c0c0",
  2470 => x"c087c401",
  2471 => x"c187c24a",
  2472 => x"2648724a",
  2473 => x"5b5e0e4f",
  2474 => x"710e5d5c",
  2475 => x"4cd4ff4b",
  2476 => x"c04866d0",
  2477 => x"ff49d678",
  2478 => x"c387d9dd",
  2479 => x"496c7cff",
  2480 => x"7199ffc3",
  2481 => x"f0c3494d",
  2482 => x"a9e0c199",
  2483 => x"c387cb05",
  2484 => x"486c7cff",
  2485 => x"66d098c3",
  2486 => x"ffc37808",
  2487 => x"494a6c7c",
  2488 => x"ffc331c8",
  2489 => x"714a6c7c",
  2490 => x"c84972b2",
  2491 => x"7cffc331",
  2492 => x"b2714a6c",
  2493 => x"31c84972",
  2494 => x"6c7cffc3",
  2495 => x"ffb2714a",
  2496 => x"e0c048d0",
  2497 => x"029b7378",
  2498 => x"7b7287c2",
  2499 => x"4d264875",
  2500 => x"4b264c26",
  2501 => x"261e4f26",
  2502 => x"5b5e0e4f",
  2503 => x"86f80e5c",
  2504 => x"a6c81e76",
  2505 => x"87fdfd49",
  2506 => x"4b7086c4",
  2507 => x"a8c4486e",
  2508 => x"87fbc203",
  2509 => x"f0c34a73",
  2510 => x"aad0c19a",
  2511 => x"c187c702",
  2512 => x"c205aae0",
  2513 => x"497387e9",
  2514 => x"c30299c8",
  2515 => x"87c6ff87",
  2516 => x"9cc34c73",
  2517 => x"c105acc2",
  2518 => x"66c487c4",
  2519 => x"7131c949",
  2520 => x"4a66c41e",
  2521 => x"c292ccc1",
  2522 => x"7249d0f7",
  2523 => x"dbcdfe81",
  2524 => x"ff49d887",
  2525 => x"c887ddda",
  2526 => x"e4c21ec0",
  2527 => x"e6fd49c8",
  2528 => x"d0ff87f1",
  2529 => x"78e0c048",
  2530 => x"1ec8e4c2",
  2531 => x"c14a66cc",
  2532 => x"f7c292cc",
  2533 => x"817249d0",
  2534 => x"87f1cbfe",
  2535 => x"acc186cc",
  2536 => x"87cbc105",
  2537 => x"fd49eec0",
  2538 => x"c487e1e3",
  2539 => x"31c94966",
  2540 => x"66c41e71",
  2541 => x"92ccc14a",
  2542 => x"49d0f7c2",
  2543 => x"ccfe8172",
  2544 => x"e4c287ca",
  2545 => x"66c81ec8",
  2546 => x"92ccc14a",
  2547 => x"49d0f7c2",
  2548 => x"c9fe8172",
  2549 => x"49d787f8",
  2550 => x"87f8d8ff",
  2551 => x"c21ec0c8",
  2552 => x"fd49c8e4",
  2553 => x"cc87e9e4",
  2554 => x"48d0ff86",
  2555 => x"f878e0c0",
  2556 => x"264c268e",
  2557 => x"1e4f264b",
  2558 => x"b7c44a71",
  2559 => x"87ce03aa",
  2560 => x"ccc14972",
  2561 => x"d0f7c291",
  2562 => x"81c8c181",
  2563 => x"4f2679c0",
  2564 => x"5c5b5e0e",
  2565 => x"86fc0e5d",
  2566 => x"d4ff4a71",
  2567 => x"d44cc04b",
  2568 => x"b7c34d66",
  2569 => x"c2c201ad",
  2570 => x"029a7287",
  2571 => x"1e87ecc0",
  2572 => x"ccc14975",
  2573 => x"d0f7c291",
  2574 => x"c8807148",
  2575 => x"66c458a6",
  2576 => x"d3c3fe49",
  2577 => x"7086c487",
  2578 => x"87d40298",
  2579 => x"c8c1496e",
  2580 => x"6e79c181",
  2581 => x"6981c849",
  2582 => x"7587c54c",
  2583 => x"87d7fe49",
  2584 => x"c848d0ff",
  2585 => x"7bdd78e1",
  2586 => x"ffc34874",
  2587 => x"747b7098",
  2588 => x"29b7c849",
  2589 => x"ffc34871",
  2590 => x"747b7098",
  2591 => x"29b7d049",
  2592 => x"ffc34871",
  2593 => x"747b7098",
  2594 => x"28b7d848",
  2595 => x"7bc07b70",
  2596 => x"7b7b7b7b",
  2597 => x"7b7b7b7b",
  2598 => x"ff7b7b7b",
  2599 => x"e0c048d0",
  2600 => x"dc1e7578",
  2601 => x"d0d6ff49",
  2602 => x"fc86c487",
  2603 => x"264d268e",
  2604 => x"264b264c",
  2605 => x"e3c21e4f",
  2606 => x"fe49bfc4",
  2607 => x"c087c3dd",
  2608 => x"004f2648",
  2609 => x"000028c8",
  2610 => x"43455053",
  2611 => x"4d555254",
  2612 => x"004d4f52",
  2613 => x"00001bbf",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
