
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"fc",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"c0",x"fc",x"c2"),
    18 => (x"48",x"d8",x"e3",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"d8",x"e3",x"c2",x"87"),
    25 => (x"d4",x"e3",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e8",x"c1",x"87",x"f7"),
    29 => (x"e3",x"c2",x"87",x"fb"),
    30 => (x"e3",x"c2",x"4d",x"d8"),
    31 => (x"ad",x"74",x"4c",x"d8"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"81",x"48",x"73",x"1e"),
    65 => (x"c5",x"02",x"a9",x"73"),
    66 => (x"05",x"53",x"12",x"87"),
    67 => (x"4f",x"26",x"87",x"f6"),
    68 => (x"71",x"1e",x"73",x"1e"),
    69 => (x"4b",x"66",x"c8",x"4a"),
    70 => (x"71",x"8b",x"c1",x"49"),
    71 => (x"87",x"cf",x"02",x"99"),
    72 => (x"d4",x"ff",x"48",x"12"),
    73 => (x"49",x"73",x"78",x"08"),
    74 => (x"99",x"71",x"8b",x"c1"),
    75 => (x"26",x"87",x"f1",x"05"),
    76 => (x"0e",x"4f",x"26",x"4b"),
    77 => (x"0e",x"5c",x"5b",x"5e"),
    78 => (x"d4",x"ff",x"4a",x"71"),
    79 => (x"4b",x"66",x"cc",x"4c"),
    80 => (x"71",x"8b",x"c1",x"49"),
    81 => (x"87",x"ce",x"02",x"99"),
    82 => (x"6c",x"7c",x"ff",x"c3"),
    83 => (x"c1",x"49",x"73",x"52"),
    84 => (x"05",x"99",x"71",x"8b"),
    85 => (x"4c",x"26",x"87",x"f2"),
    86 => (x"4f",x"26",x"4b",x"26"),
    87 => (x"ff",x"1e",x"73",x"1e"),
    88 => (x"ff",x"c3",x"4b",x"d4"),
    89 => (x"c3",x"4a",x"6b",x"7b"),
    90 => (x"49",x"6b",x"7b",x"ff"),
    91 => (x"b1",x"72",x"32",x"c8"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"71",x"31",x"c8",x"4a"),
    94 => (x"7b",x"ff",x"c3",x"b2"),
    95 => (x"32",x"c8",x"49",x"6b"),
    96 => (x"48",x"71",x"b1",x"72"),
    97 => (x"4f",x"26",x"4b",x"26"),
    98 => (x"5c",x"5b",x"5e",x"0e"),
    99 => (x"4d",x"71",x"0e",x"5d"),
   100 => (x"75",x"4c",x"d4",x"ff"),
   101 => (x"98",x"ff",x"c3",x"48"),
   102 => (x"e3",x"c2",x"7c",x"70"),
   103 => (x"c8",x"05",x"bf",x"d8"),
   104 => (x"48",x"66",x"d0",x"87"),
   105 => (x"a6",x"d4",x"30",x"c9"),
   106 => (x"49",x"66",x"d0",x"58"),
   107 => (x"48",x"71",x"29",x"d8"),
   108 => (x"70",x"98",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"48",x"71",x"29",x"d0"),
   111 => (x"70",x"98",x"ff",x"c3"),
   112 => (x"49",x"66",x"d0",x"7c"),
   113 => (x"48",x"71",x"29",x"c8"),
   114 => (x"70",x"98",x"ff",x"c3"),
   115 => (x"48",x"66",x"d0",x"7c"),
   116 => (x"70",x"98",x"ff",x"c3"),
   117 => (x"d0",x"49",x"75",x"7c"),
   118 => (x"c3",x"48",x"71",x"29"),
   119 => (x"7c",x"70",x"98",x"ff"),
   120 => (x"f0",x"c9",x"4b",x"6c"),
   121 => (x"ff",x"c3",x"4a",x"ff"),
   122 => (x"87",x"cf",x"05",x"ab"),
   123 => (x"6c",x"7c",x"71",x"49"),
   124 => (x"02",x"8a",x"c1",x"4b"),
   125 => (x"ab",x"71",x"87",x"c5"),
   126 => (x"73",x"87",x"f2",x"02"),
   127 => (x"26",x"4d",x"26",x"48"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"49",x"c0",x"1e",x"4f"),
   130 => (x"c3",x"48",x"d4",x"ff"),
   131 => (x"81",x"c1",x"78",x"ff"),
   132 => (x"a9",x"b7",x"c8",x"c3"),
   133 => (x"26",x"87",x"f1",x"04"),
   134 => (x"5b",x"5e",x"0e",x"4f"),
   135 => (x"c0",x"0e",x"5d",x"5c"),
   136 => (x"f7",x"c1",x"f0",x"ff"),
   137 => (x"c0",x"c0",x"c1",x"4d"),
   138 => (x"4b",x"c0",x"c0",x"c0"),
   139 => (x"c4",x"87",x"d6",x"ff"),
   140 => (x"c0",x"4c",x"df",x"f8"),
   141 => (x"fd",x"49",x"75",x"1e"),
   142 => (x"86",x"c4",x"87",x"ce"),
   143 => (x"c0",x"05",x"a8",x"c1"),
   144 => (x"d4",x"ff",x"87",x"e5"),
   145 => (x"78",x"ff",x"c3",x"48"),
   146 => (x"e1",x"c0",x"1e",x"73"),
   147 => (x"49",x"e9",x"c1",x"f0"),
   148 => (x"c4",x"87",x"f5",x"fc"),
   149 => (x"05",x"98",x"70",x"86"),
   150 => (x"d4",x"ff",x"87",x"ca"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"87",x"cb",x"48",x"c1"),
   153 => (x"c1",x"87",x"de",x"fe"),
   154 => (x"c6",x"ff",x"05",x"8c"),
   155 => (x"26",x"48",x"c0",x"87"),
   156 => (x"26",x"4c",x"26",x"4d"),
   157 => (x"0e",x"4f",x"26",x"4b"),
   158 => (x"0e",x"5c",x"5b",x"5e"),
   159 => (x"c1",x"f0",x"ff",x"c0"),
   160 => (x"d4",x"ff",x"4c",x"c1"),
   161 => (x"78",x"ff",x"c3",x"48"),
   162 => (x"f8",x"49",x"fc",x"ca"),
   163 => (x"4b",x"d3",x"87",x"d9"),
   164 => (x"49",x"74",x"1e",x"c0"),
   165 => (x"c4",x"87",x"f1",x"fb"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"d4",x"ff",x"87",x"ca"),
   168 => (x"78",x"ff",x"c3",x"48"),
   169 => (x"87",x"cb",x"48",x"c1"),
   170 => (x"c1",x"87",x"da",x"fd"),
   171 => (x"df",x"ff",x"05",x"8b"),
   172 => (x"26",x"48",x"c0",x"87"),
   173 => (x"26",x"4b",x"26",x"4c"),
   174 => (x"00",x"00",x"00",x"4f"),
   175 => (x"00",x"44",x"4d",x"43"),
   176 => (x"43",x"48",x"44",x"53"),
   177 => (x"69",x"61",x"66",x"20"),
   178 => (x"00",x"0a",x"21",x"6c"),
   179 => (x"52",x"52",x"45",x"49"),
   180 => (x"00",x"00",x"00",x"00"),
   181 => (x"00",x"49",x"50",x"53"),
   182 => (x"74",x"69",x"72",x"57"),
   183 => (x"61",x"66",x"20",x"65"),
   184 => (x"64",x"65",x"6c",x"69"),
   185 => (x"5e",x"0e",x"00",x"0a"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"d0",x"fc",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"c7",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"ec",x"fd"),
   195 => (x"87",x"e8",x"c1",x"48"),
   196 => (x"70",x"87",x"c9",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fd",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"d5"),
   201 => (x"75",x"87",x"d1",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"ea",x"fb"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"c8",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"db",x"48",x"c1",x"87"),
   215 => (x"d7",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"c0",x"cb",x"87",x"ca"),
   218 => (x"87",x"fb",x"f4",x"49"),
   219 => (x"87",x"c8",x"48",x"c0"),
   220 => (x"fe",x"05",x"8c",x"c1"),
   221 => (x"48",x"c0",x"87",x"f6"),
   222 => (x"4c",x"26",x"4d",x"26"),
   223 => (x"4f",x"26",x"4b",x"26"),
   224 => (x"5c",x"5b",x"5e",x"0e"),
   225 => (x"d0",x"ff",x"0e",x"5d"),
   226 => (x"d0",x"e5",x"c0",x"4d"),
   227 => (x"c2",x"4c",x"c0",x"c1"),
   228 => (x"c1",x"48",x"d8",x"e3"),
   229 => (x"49",x"d4",x"cb",x"78"),
   230 => (x"c7",x"87",x"cc",x"f4"),
   231 => (x"f9",x"7d",x"c2",x"4b"),
   232 => (x"7d",x"c3",x"87",x"e3"),
   233 => (x"49",x"74",x"1e",x"c0"),
   234 => (x"c4",x"87",x"dd",x"f7"),
   235 => (x"05",x"a8",x"c1",x"86"),
   236 => (x"c2",x"4b",x"87",x"c1"),
   237 => (x"87",x"cb",x"05",x"ab"),
   238 => (x"f3",x"49",x"cc",x"cb"),
   239 => (x"48",x"c0",x"87",x"e9"),
   240 => (x"c1",x"87",x"f6",x"c0"),
   241 => (x"d4",x"ff",x"05",x"8b"),
   242 => (x"87",x"da",x"fc",x"87"),
   243 => (x"58",x"dc",x"e3",x"c2"),
   244 => (x"cd",x"05",x"98",x"70"),
   245 => (x"c0",x"1e",x"c1",x"87"),
   246 => (x"d0",x"c1",x"f0",x"ff"),
   247 => (x"87",x"e8",x"f6",x"49"),
   248 => (x"d4",x"ff",x"86",x"c4"),
   249 => (x"78",x"ff",x"c3",x"48"),
   250 => (x"c2",x"87",x"ee",x"c4"),
   251 => (x"c2",x"58",x"e0",x"e3"),
   252 => (x"48",x"d4",x"ff",x"7d"),
   253 => (x"c1",x"78",x"ff",x"c3"),
   254 => (x"26",x"4d",x"26",x"48"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"71",x"0e",x"5d",x"5c"),
   258 => (x"4c",x"ff",x"c3",x"4d"),
   259 => (x"74",x"4b",x"d4",x"ff"),
   260 => (x"48",x"d0",x"ff",x"7b"),
   261 => (x"74",x"78",x"c3",x"c4"),
   262 => (x"c0",x"1e",x"75",x"7b"),
   263 => (x"d8",x"c1",x"f0",x"ff"),
   264 => (x"87",x"e4",x"f5",x"49"),
   265 => (x"98",x"70",x"86",x"c4"),
   266 => (x"cb",x"87",x"cb",x"02"),
   267 => (x"f6",x"f1",x"49",x"d8"),
   268 => (x"c0",x"48",x"c1",x"87"),
   269 => (x"7b",x"74",x"87",x"ee"),
   270 => (x"c8",x"7b",x"fe",x"c3"),
   271 => (x"66",x"d4",x"1e",x"c0"),
   272 => (x"87",x"cc",x"f3",x"49"),
   273 => (x"7b",x"74",x"86",x"c4"),
   274 => (x"7b",x"74",x"7b",x"74"),
   275 => (x"4a",x"e0",x"da",x"d8"),
   276 => (x"05",x"6b",x"7b",x"74"),
   277 => (x"8a",x"c1",x"87",x"c5"),
   278 => (x"74",x"87",x"f5",x"05"),
   279 => (x"48",x"d0",x"ff",x"7b"),
   280 => (x"48",x"c0",x"78",x"c2"),
   281 => (x"4c",x"26",x"4d",x"26"),
   282 => (x"4f",x"26",x"4b",x"26"),
   283 => (x"5c",x"5b",x"5e",x"0e"),
   284 => (x"86",x"fc",x"0e",x"5d"),
   285 => (x"d4",x"ff",x"4b",x"71"),
   286 => (x"c5",x"7e",x"c0",x"4c"),
   287 => (x"4a",x"df",x"cd",x"ee"),
   288 => (x"6c",x"7c",x"ff",x"c3"),
   289 => (x"a8",x"fe",x"c3",x"48"),
   290 => (x"87",x"f8",x"c0",x"05"),
   291 => (x"9b",x"73",x"4d",x"74"),
   292 => (x"d4",x"87",x"cc",x"02"),
   293 => (x"49",x"73",x"1e",x"66"),
   294 => (x"c4",x"87",x"d8",x"f2"),
   295 => (x"ff",x"87",x"d4",x"86"),
   296 => (x"d1",x"c4",x"48",x"d0"),
   297 => (x"4a",x"66",x"d4",x"78"),
   298 => (x"c1",x"7d",x"ff",x"c3"),
   299 => (x"87",x"f8",x"05",x"8a"),
   300 => (x"c3",x"5a",x"a6",x"d8"),
   301 => (x"73",x"7c",x"7c",x"ff"),
   302 => (x"87",x"c5",x"05",x"9b"),
   303 => (x"d0",x"48",x"d0",x"ff"),
   304 => (x"7e",x"4a",x"c1",x"78"),
   305 => (x"fe",x"05",x"8a",x"c1"),
   306 => (x"48",x"6e",x"87",x"f6"),
   307 => (x"4d",x"26",x"8e",x"fc"),
   308 => (x"4b",x"26",x"4c",x"26"),
   309 => (x"73",x"1e",x"4f",x"26"),
   310 => (x"c0",x"4a",x"71",x"1e"),
   311 => (x"48",x"d4",x"ff",x"4b"),
   312 => (x"ff",x"78",x"ff",x"c3"),
   313 => (x"c3",x"c4",x"48",x"d0"),
   314 => (x"48",x"d4",x"ff",x"78"),
   315 => (x"72",x"78",x"ff",x"c3"),
   316 => (x"f0",x"ff",x"c0",x"1e"),
   317 => (x"f2",x"49",x"d1",x"c1"),
   318 => (x"86",x"c4",x"87",x"ce"),
   319 => (x"d2",x"05",x"98",x"70"),
   320 => (x"1e",x"c0",x"c8",x"87"),
   321 => (x"fd",x"49",x"66",x"cc"),
   322 => (x"86",x"c4",x"87",x"e2"),
   323 => (x"d0",x"ff",x"4b",x"70"),
   324 => (x"73",x"78",x"c2",x"48"),
   325 => (x"26",x"4b",x"26",x"48"),
   326 => (x"5b",x"5e",x"0e",x"4f"),
   327 => (x"c0",x"0e",x"5d",x"5c"),
   328 => (x"f0",x"ff",x"c0",x"1e"),
   329 => (x"f1",x"49",x"c9",x"c1"),
   330 => (x"1e",x"d2",x"87",x"de"),
   331 => (x"49",x"e8",x"e3",x"c2"),
   332 => (x"c8",x"87",x"f9",x"fc"),
   333 => (x"c1",x"4c",x"c0",x"86"),
   334 => (x"ac",x"b7",x"d2",x"84"),
   335 => (x"c2",x"87",x"f8",x"04"),
   336 => (x"bf",x"97",x"e8",x"e3"),
   337 => (x"99",x"c0",x"c3",x"49"),
   338 => (x"05",x"a9",x"c0",x"c1"),
   339 => (x"c2",x"87",x"e7",x"c0"),
   340 => (x"bf",x"97",x"ef",x"e3"),
   341 => (x"c2",x"31",x"d0",x"49"),
   342 => (x"bf",x"97",x"f0",x"e3"),
   343 => (x"72",x"32",x"c8",x"4a"),
   344 => (x"f1",x"e3",x"c2",x"b1"),
   345 => (x"b1",x"4a",x"bf",x"97"),
   346 => (x"ff",x"cf",x"4c",x"71"),
   347 => (x"c1",x"9c",x"ff",x"ff"),
   348 => (x"c1",x"34",x"ca",x"84"),
   349 => (x"e3",x"c2",x"87",x"e7"),
   350 => (x"49",x"bf",x"97",x"f1"),
   351 => (x"99",x"c6",x"31",x"c1"),
   352 => (x"97",x"f2",x"e3",x"c2"),
   353 => (x"b7",x"c7",x"4a",x"bf"),
   354 => (x"c2",x"b1",x"72",x"2a"),
   355 => (x"bf",x"97",x"ed",x"e3"),
   356 => (x"9d",x"cf",x"4d",x"4a"),
   357 => (x"97",x"ee",x"e3",x"c2"),
   358 => (x"9a",x"c3",x"4a",x"bf"),
   359 => (x"e3",x"c2",x"32",x"ca"),
   360 => (x"4b",x"bf",x"97",x"ef"),
   361 => (x"b2",x"73",x"33",x"c2"),
   362 => (x"97",x"f0",x"e3",x"c2"),
   363 => (x"c0",x"c3",x"4b",x"bf"),
   364 => (x"2b",x"b7",x"c6",x"9b"),
   365 => (x"81",x"c2",x"b2",x"73"),
   366 => (x"30",x"71",x"48",x"c1"),
   367 => (x"48",x"c1",x"49",x"70"),
   368 => (x"4d",x"70",x"30",x"75"),
   369 => (x"84",x"c1",x"4c",x"72"),
   370 => (x"c0",x"c8",x"94",x"71"),
   371 => (x"cc",x"06",x"ad",x"b7"),
   372 => (x"b7",x"34",x"c1",x"87"),
   373 => (x"b7",x"c0",x"c8",x"2d"),
   374 => (x"f4",x"ff",x"01",x"ad"),
   375 => (x"26",x"48",x"74",x"87"),
   376 => (x"26",x"4c",x"26",x"4d"),
   377 => (x"0e",x"4f",x"26",x"4b"),
   378 => (x"5d",x"5c",x"5b",x"5e"),
   379 => (x"c2",x"86",x"fc",x"0e"),
   380 => (x"c0",x"48",x"d0",x"ec"),
   381 => (x"c8",x"e4",x"c2",x"78"),
   382 => (x"fb",x"49",x"c0",x"1e"),
   383 => (x"86",x"c4",x"87",x"d8"),
   384 => (x"c5",x"05",x"98",x"70"),
   385 => (x"c9",x"48",x"c0",x"87"),
   386 => (x"4d",x"c0",x"87",x"d2"),
   387 => (x"48",x"cc",x"f1",x"c2"),
   388 => (x"e4",x"c2",x"78",x"c1"),
   389 => (x"e1",x"c0",x"4a",x"fe"),
   390 => (x"4b",x"c8",x"49",x"f4"),
   391 => (x"70",x"87",x"c7",x"eb"),
   392 => (x"87",x"c6",x"05",x"98"),
   393 => (x"48",x"cc",x"f1",x"c2"),
   394 => (x"e5",x"c2",x"78",x"c0"),
   395 => (x"e2",x"c0",x"4a",x"da"),
   396 => (x"4b",x"c8",x"49",x"c0"),
   397 => (x"70",x"87",x"ef",x"ea"),
   398 => (x"87",x"c6",x"05",x"98"),
   399 => (x"48",x"cc",x"f1",x"c2"),
   400 => (x"f1",x"c2",x"78",x"c0"),
   401 => (x"c0",x"02",x"bf",x"cc"),
   402 => (x"eb",x"c2",x"87",x"fd"),
   403 => (x"c2",x"4d",x"bf",x"ce"),
   404 => (x"bf",x"9f",x"c6",x"ec"),
   405 => (x"d6",x"c5",x"48",x"7e"),
   406 => (x"c7",x"05",x"a8",x"ea"),
   407 => (x"ce",x"eb",x"c2",x"87"),
   408 => (x"87",x"ce",x"4d",x"bf"),
   409 => (x"e9",x"ca",x"48",x"6e"),
   410 => (x"c5",x"02",x"a8",x"d5"),
   411 => (x"c7",x"48",x"c0",x"87"),
   412 => (x"e4",x"c2",x"87",x"ea"),
   413 => (x"49",x"75",x"1e",x"c8"),
   414 => (x"c4",x"87",x"db",x"f9"),
   415 => (x"05",x"98",x"70",x"86"),
   416 => (x"48",x"c0",x"87",x"c5"),
   417 => (x"c2",x"87",x"d5",x"c7"),
   418 => (x"c0",x"4a",x"da",x"e5"),
   419 => (x"c8",x"49",x"cc",x"e2"),
   420 => (x"87",x"d2",x"e9",x"4b"),
   421 => (x"c8",x"05",x"98",x"70"),
   422 => (x"d0",x"ec",x"c2",x"87"),
   423 => (x"d8",x"78",x"c1",x"48"),
   424 => (x"fe",x"e4",x"c2",x"87"),
   425 => (x"d8",x"e2",x"c0",x"4a"),
   426 => (x"e8",x"4b",x"c8",x"49"),
   427 => (x"98",x"70",x"87",x"f8"),
   428 => (x"87",x"c5",x"c0",x"02"),
   429 => (x"e3",x"c6",x"48",x"c0"),
   430 => (x"c6",x"ec",x"c2",x"87"),
   431 => (x"c1",x"49",x"bf",x"97"),
   432 => (x"c0",x"05",x"a9",x"d5"),
   433 => (x"ec",x"c2",x"87",x"cd"),
   434 => (x"49",x"bf",x"97",x"c7"),
   435 => (x"02",x"a9",x"ea",x"c2"),
   436 => (x"c0",x"87",x"c5",x"c0"),
   437 => (x"87",x"c4",x"c6",x"48"),
   438 => (x"97",x"c8",x"e4",x"c2"),
   439 => (x"c3",x"48",x"7e",x"bf"),
   440 => (x"c0",x"02",x"a8",x"e9"),
   441 => (x"48",x"6e",x"87",x"ce"),
   442 => (x"02",x"a8",x"eb",x"c3"),
   443 => (x"c0",x"87",x"c5",x"c0"),
   444 => (x"87",x"e8",x"c5",x"48"),
   445 => (x"97",x"d3",x"e4",x"c2"),
   446 => (x"05",x"99",x"49",x"bf"),
   447 => (x"c2",x"87",x"cc",x"c0"),
   448 => (x"bf",x"97",x"d4",x"e4"),
   449 => (x"02",x"a9",x"c2",x"49"),
   450 => (x"c0",x"87",x"c5",x"c0"),
   451 => (x"87",x"cc",x"c5",x"48"),
   452 => (x"97",x"d5",x"e4",x"c2"),
   453 => (x"ec",x"c2",x"48",x"bf"),
   454 => (x"4c",x"70",x"58",x"cc"),
   455 => (x"c2",x"88",x"c1",x"48"),
   456 => (x"c2",x"58",x"d0",x"ec"),
   457 => (x"bf",x"97",x"d6",x"e4"),
   458 => (x"c2",x"81",x"75",x"49"),
   459 => (x"bf",x"97",x"d7",x"e4"),
   460 => (x"72",x"32",x"c8",x"4a"),
   461 => (x"f0",x"c2",x"7e",x"a1"),
   462 => (x"78",x"6e",x"48",x"e8"),
   463 => (x"97",x"d8",x"e4",x"c2"),
   464 => (x"f1",x"c2",x"48",x"bf"),
   465 => (x"ec",x"c2",x"58",x"c0"),
   466 => (x"c2",x"02",x"bf",x"d0"),
   467 => (x"e5",x"c2",x"87",x"d3"),
   468 => (x"e1",x"c0",x"4a",x"da"),
   469 => (x"4b",x"c8",x"49",x"e8"),
   470 => (x"70",x"87",x"cb",x"e6"),
   471 => (x"c5",x"c0",x"02",x"98"),
   472 => (x"c3",x"48",x"c0",x"87"),
   473 => (x"ec",x"c2",x"87",x"f6"),
   474 => (x"c2",x"4c",x"bf",x"c8"),
   475 => (x"c2",x"5c",x"fc",x"f0"),
   476 => (x"bf",x"97",x"ed",x"e4"),
   477 => (x"c2",x"31",x"c8",x"49"),
   478 => (x"bf",x"97",x"ec",x"e4"),
   479 => (x"c2",x"49",x"a1",x"4a"),
   480 => (x"bf",x"97",x"ee",x"e4"),
   481 => (x"72",x"32",x"d0",x"4a"),
   482 => (x"e4",x"c2",x"49",x"a1"),
   483 => (x"4a",x"bf",x"97",x"ef"),
   484 => (x"a1",x"72",x"32",x"d8"),
   485 => (x"c4",x"f1",x"c2",x"49"),
   486 => (x"fc",x"f0",x"c2",x"59"),
   487 => (x"f0",x"c2",x"91",x"bf"),
   488 => (x"c2",x"81",x"bf",x"e8"),
   489 => (x"c2",x"59",x"f0",x"f0"),
   490 => (x"bf",x"97",x"f5",x"e4"),
   491 => (x"c2",x"32",x"c8",x"4a"),
   492 => (x"bf",x"97",x"f4",x"e4"),
   493 => (x"c2",x"4a",x"a2",x"4b"),
   494 => (x"bf",x"97",x"f6",x"e4"),
   495 => (x"73",x"33",x"d0",x"4b"),
   496 => (x"e4",x"c2",x"4a",x"a2"),
   497 => (x"4b",x"bf",x"97",x"f7"),
   498 => (x"33",x"d8",x"9b",x"cf"),
   499 => (x"c2",x"4a",x"a2",x"73"),
   500 => (x"c2",x"5a",x"f4",x"f0"),
   501 => (x"c2",x"92",x"74",x"8a"),
   502 => (x"72",x"48",x"f4",x"f0"),
   503 => (x"c7",x"c1",x"78",x"a1"),
   504 => (x"da",x"e4",x"c2",x"87"),
   505 => (x"c8",x"49",x"bf",x"97"),
   506 => (x"d9",x"e4",x"c2",x"31"),
   507 => (x"a1",x"4a",x"bf",x"97"),
   508 => (x"c7",x"31",x"c5",x"49"),
   509 => (x"29",x"c9",x"81",x"ff"),
   510 => (x"59",x"fc",x"f0",x"c2"),
   511 => (x"97",x"df",x"e4",x"c2"),
   512 => (x"32",x"c8",x"4a",x"bf"),
   513 => (x"97",x"de",x"e4",x"c2"),
   514 => (x"4a",x"a2",x"4b",x"bf"),
   515 => (x"5a",x"c4",x"f1",x"c2"),
   516 => (x"bf",x"fc",x"f0",x"c2"),
   517 => (x"c2",x"82",x"6e",x"92"),
   518 => (x"c2",x"5a",x"f8",x"f0"),
   519 => (x"c0",x"48",x"f0",x"f0"),
   520 => (x"ec",x"f0",x"c2",x"78"),
   521 => (x"78",x"a1",x"72",x"48"),
   522 => (x"48",x"c4",x"f1",x"c2"),
   523 => (x"bf",x"f0",x"f0",x"c2"),
   524 => (x"c8",x"f1",x"c2",x"78"),
   525 => (x"f4",x"f0",x"c2",x"48"),
   526 => (x"ec",x"c2",x"78",x"bf"),
   527 => (x"c0",x"02",x"bf",x"d0"),
   528 => (x"48",x"74",x"87",x"c9"),
   529 => (x"7e",x"70",x"30",x"c4"),
   530 => (x"c2",x"87",x"c9",x"c0"),
   531 => (x"48",x"bf",x"f8",x"f0"),
   532 => (x"7e",x"70",x"30",x"c4"),
   533 => (x"48",x"d4",x"ec",x"c2"),
   534 => (x"48",x"c1",x"78",x"6e"),
   535 => (x"4d",x"26",x"8e",x"fc"),
   536 => (x"4b",x"26",x"4c",x"26"),
   537 => (x"00",x"00",x"4f",x"26"),
   538 => (x"33",x"54",x"41",x"46"),
   539 => (x"20",x"20",x"20",x"32"),
   540 => (x"00",x"00",x"00",x"00"),
   541 => (x"31",x"54",x"41",x"46"),
   542 => (x"20",x"20",x"20",x"36"),
   543 => (x"00",x"00",x"00",x"00"),
   544 => (x"33",x"54",x"41",x"46"),
   545 => (x"20",x"20",x"20",x"32"),
   546 => (x"00",x"00",x"00",x"00"),
   547 => (x"33",x"54",x"41",x"46"),
   548 => (x"20",x"20",x"20",x"32"),
   549 => (x"00",x"00",x"00",x"00"),
   550 => (x"31",x"54",x"41",x"46"),
   551 => (x"20",x"20",x"20",x"36"),
   552 => (x"5b",x"5e",x"0e",x"00"),
   553 => (x"71",x"0e",x"5d",x"5c"),
   554 => (x"d0",x"ec",x"c2",x"4a"),
   555 => (x"87",x"cb",x"02",x"bf"),
   556 => (x"2b",x"c7",x"4b",x"72"),
   557 => (x"ff",x"c1",x"4d",x"72"),
   558 => (x"72",x"87",x"c9",x"9d"),
   559 => (x"72",x"2b",x"c8",x"4b"),
   560 => (x"9d",x"ff",x"c3",x"4d"),
   561 => (x"bf",x"e8",x"f0",x"c2"),
   562 => (x"e8",x"f9",x"c0",x"83"),
   563 => (x"d9",x"02",x"ab",x"bf"),
   564 => (x"ec",x"f9",x"c0",x"87"),
   565 => (x"c8",x"e4",x"c2",x"5b"),
   566 => (x"ef",x"49",x"73",x"1e"),
   567 => (x"86",x"c4",x"87",x"f8"),
   568 => (x"c5",x"05",x"98",x"70"),
   569 => (x"c0",x"48",x"c0",x"87"),
   570 => (x"ec",x"c2",x"87",x"e6"),
   571 => (x"d2",x"02",x"bf",x"d0"),
   572 => (x"c4",x"49",x"75",x"87"),
   573 => (x"c8",x"e4",x"c2",x"91"),
   574 => (x"cf",x"4c",x"69",x"81"),
   575 => (x"ff",x"ff",x"ff",x"ff"),
   576 => (x"75",x"87",x"cb",x"9c"),
   577 => (x"c2",x"91",x"c2",x"49"),
   578 => (x"9f",x"81",x"c8",x"e4"),
   579 => (x"48",x"74",x"4c",x"69"),
   580 => (x"4c",x"26",x"4d",x"26"),
   581 => (x"4f",x"26",x"4b",x"26"),
   582 => (x"5c",x"5b",x"5e",x"0e"),
   583 => (x"86",x"f4",x"0e",x"5d"),
   584 => (x"c4",x"59",x"a6",x"c8"),
   585 => (x"80",x"c8",x"48",x"66"),
   586 => (x"c0",x"48",x"7e",x"70"),
   587 => (x"49",x"c1",x"1e",x"78"),
   588 => (x"87",x"f9",x"cc",x"49"),
   589 => (x"4c",x"70",x"86",x"c4"),
   590 => (x"fc",x"c0",x"02",x"9c"),
   591 => (x"d8",x"ec",x"c2",x"87"),
   592 => (x"49",x"66",x"dc",x"4a"),
   593 => (x"87",x"c3",x"de",x"ff"),
   594 => (x"c0",x"02",x"98",x"70"),
   595 => (x"4a",x"74",x"87",x"eb"),
   596 => (x"cb",x"49",x"66",x"dc"),
   597 => (x"cd",x"de",x"ff",x"4b"),
   598 => (x"02",x"98",x"70",x"87"),
   599 => (x"1e",x"c0",x"87",x"db"),
   600 => (x"c4",x"02",x"9c",x"74"),
   601 => (x"c2",x"4d",x"c0",x"87"),
   602 => (x"75",x"4d",x"c1",x"87"),
   603 => (x"87",x"fd",x"cb",x"49"),
   604 => (x"4c",x"70",x"86",x"c4"),
   605 => (x"c4",x"ff",x"05",x"9c"),
   606 => (x"02",x"9c",x"74",x"87"),
   607 => (x"dc",x"87",x"f4",x"c1"),
   608 => (x"48",x"6e",x"49",x"a4"),
   609 => (x"a4",x"da",x"78",x"69"),
   610 => (x"4d",x"66",x"c4",x"49"),
   611 => (x"69",x"9f",x"85",x"c4"),
   612 => (x"d0",x"ec",x"c2",x"7d"),
   613 => (x"87",x"d2",x"02",x"bf"),
   614 => (x"9f",x"49",x"a4",x"d4"),
   615 => (x"ff",x"c0",x"49",x"69"),
   616 => (x"48",x"71",x"99",x"ff"),
   617 => (x"7e",x"70",x"30",x"d0"),
   618 => (x"7e",x"c0",x"87",x"c2"),
   619 => (x"6d",x"48",x"49",x"6e"),
   620 => (x"c4",x"7d",x"70",x"80"),
   621 => (x"78",x"c0",x"48",x"66"),
   622 => (x"cc",x"49",x"66",x"c4"),
   623 => (x"c4",x"79",x"6d",x"81"),
   624 => (x"81",x"d0",x"49",x"66"),
   625 => (x"a6",x"c8",x"79",x"c0"),
   626 => (x"c8",x"78",x"c0",x"48"),
   627 => (x"66",x"c4",x"4c",x"66"),
   628 => (x"74",x"82",x"d4",x"4a"),
   629 => (x"72",x"91",x"c8",x"49"),
   630 => (x"41",x"c0",x"49",x"a1"),
   631 => (x"84",x"c1",x"79",x"6d"),
   632 => (x"04",x"ac",x"b7",x"c6"),
   633 => (x"c4",x"87",x"e7",x"ff"),
   634 => (x"c4",x"c1",x"49",x"66"),
   635 => (x"c1",x"79",x"c0",x"81"),
   636 => (x"c0",x"87",x"c2",x"48"),
   637 => (x"26",x"8e",x"f4",x"48"),
   638 => (x"26",x"4c",x"26",x"4d"),
   639 => (x"0e",x"4f",x"26",x"4b"),
   640 => (x"5d",x"5c",x"5b",x"5e"),
   641 => (x"d0",x"4c",x"71",x"0e"),
   642 => (x"6c",x"4a",x"4d",x"66"),
   643 => (x"4d",x"a1",x"72",x"49"),
   644 => (x"cc",x"ec",x"c2",x"b9"),
   645 => (x"ba",x"ff",x"4a",x"bf"),
   646 => (x"99",x"71",x"99",x"72"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"6b",x"4b",x"a4",x"c4"),
   649 => (x"87",x"f9",x"f9",x"49"),
   650 => (x"ec",x"c2",x"7b",x"70"),
   651 => (x"6c",x"49",x"bf",x"c8"),
   652 => (x"75",x"7c",x"71",x"81"),
   653 => (x"cc",x"ec",x"c2",x"b9"),
   654 => (x"ba",x"ff",x"4a",x"bf"),
   655 => (x"99",x"71",x"99",x"72"),
   656 => (x"87",x"dc",x"ff",x"05"),
   657 => (x"4d",x"26",x"7c",x"75"),
   658 => (x"4b",x"26",x"4c",x"26"),
   659 => (x"73",x"1e",x"4f",x"26"),
   660 => (x"c2",x"4b",x"71",x"1e"),
   661 => (x"49",x"bf",x"ec",x"f0"),
   662 => (x"6a",x"4a",x"a3",x"c4"),
   663 => (x"c2",x"8a",x"c2",x"4a"),
   664 => (x"92",x"bf",x"c8",x"ec"),
   665 => (x"c2",x"49",x"a1",x"72"),
   666 => (x"4a",x"bf",x"cc",x"ec"),
   667 => (x"a1",x"72",x"9a",x"6b"),
   668 => (x"ec",x"f9",x"c0",x"49"),
   669 => (x"1e",x"66",x"c8",x"59"),
   670 => (x"87",x"da",x"e9",x"71"),
   671 => (x"98",x"70",x"86",x"c4"),
   672 => (x"c0",x"87",x"c4",x"05"),
   673 => (x"c1",x"87",x"c2",x"48"),
   674 => (x"26",x"4b",x"26",x"48"),
   675 => (x"1e",x"73",x"1e",x"4f"),
   676 => (x"f0",x"c2",x"4b",x"71"),
   677 => (x"c4",x"49",x"bf",x"ec"),
   678 => (x"4a",x"6a",x"4a",x"a3"),
   679 => (x"ec",x"c2",x"8a",x"c2"),
   680 => (x"72",x"92",x"bf",x"c8"),
   681 => (x"ec",x"c2",x"49",x"a1"),
   682 => (x"6b",x"4a",x"bf",x"cc"),
   683 => (x"49",x"a1",x"72",x"9a"),
   684 => (x"59",x"ec",x"f9",x"c0"),
   685 => (x"71",x"1e",x"66",x"c8"),
   686 => (x"c4",x"87",x"c6",x"e5"),
   687 => (x"05",x"98",x"70",x"86"),
   688 => (x"48",x"c0",x"87",x"c4"),
   689 => (x"48",x"c1",x"87",x"c2"),
   690 => (x"4f",x"26",x"4b",x"26"),
   691 => (x"5c",x"5b",x"5e",x"0e"),
   692 => (x"86",x"e0",x"0e",x"5d"),
   693 => (x"f0",x"c0",x"4b",x"71"),
   694 => (x"29",x"c9",x"49",x"66"),
   695 => (x"c2",x"59",x"a6",x"c8"),
   696 => (x"49",x"bf",x"cc",x"ec"),
   697 => (x"4a",x"71",x"b9",x"ff"),
   698 => (x"d8",x"9a",x"66",x"c4"),
   699 => (x"99",x"6b",x"5a",x"a6"),
   700 => (x"c4",x"59",x"a6",x"d0"),
   701 => (x"a6",x"d0",x"7e",x"a3"),
   702 => (x"78",x"bf",x"6e",x"48"),
   703 => (x"cc",x"48",x"66",x"d4"),
   704 => (x"c6",x"05",x"a8",x"66"),
   705 => (x"7b",x"66",x"c4",x"87"),
   706 => (x"d8",x"87",x"c1",x"c3"),
   707 => (x"ff",x"c1",x"48",x"a6"),
   708 => (x"ff",x"ff",x"ff",x"ff"),
   709 => (x"ff",x"80",x"c4",x"78"),
   710 => (x"c8",x"4c",x"c0",x"78"),
   711 => (x"a3",x"d4",x"48",x"a6"),
   712 => (x"c8",x"49",x"74",x"78"),
   713 => (x"81",x"66",x"c8",x"91"),
   714 => (x"4d",x"4a",x"66",x"d4"),
   715 => (x"b7",x"c0",x"8d",x"69"),
   716 => (x"87",x"ce",x"04",x"ad"),
   717 => (x"ad",x"b7",x"66",x"d8"),
   718 => (x"c0",x"87",x"c7",x"03"),
   719 => (x"dc",x"5c",x"a6",x"e0"),
   720 => (x"84",x"c1",x"5d",x"a6"),
   721 => (x"04",x"ac",x"b7",x"c6"),
   722 => (x"dc",x"87",x"d0",x"ff"),
   723 => (x"b7",x"c0",x"48",x"66"),
   724 => (x"87",x"d0",x"04",x"a8"),
   725 => (x"c8",x"49",x"66",x"dc"),
   726 => (x"81",x"66",x"c8",x"91"),
   727 => (x"48",x"6e",x"7b",x"21"),
   728 => (x"87",x"c9",x"78",x"69"),
   729 => (x"a3",x"cc",x"7b",x"c0"),
   730 => (x"69",x"48",x"6e",x"49"),
   731 => (x"48",x"66",x"c4",x"78"),
   732 => (x"a6",x"c8",x"88",x"6b"),
   733 => (x"c8",x"ec",x"c2",x"58"),
   734 => (x"90",x"c8",x"48",x"bf"),
   735 => (x"66",x"c4",x"7e",x"70"),
   736 => (x"01",x"a8",x"6e",x"48"),
   737 => (x"66",x"c4",x"87",x"c9"),
   738 => (x"03",x"a8",x"6e",x"48"),
   739 => (x"c1",x"87",x"f3",x"c0"),
   740 => (x"6a",x"4a",x"a3",x"c4"),
   741 => (x"c8",x"91",x"c8",x"49"),
   742 => (x"66",x"cc",x"81",x"66"),
   743 => (x"c8",x"49",x"6a",x"79"),
   744 => (x"81",x"66",x"c8",x"91"),
   745 => (x"66",x"d0",x"81",x"c4"),
   746 => (x"48",x"7e",x"6a",x"79"),
   747 => (x"c7",x"05",x"a8",x"c5"),
   748 => (x"48",x"a6",x"c8",x"87"),
   749 => (x"87",x"c7",x"78",x"c0"),
   750 => (x"80",x"c1",x"48",x"6e"),
   751 => (x"c8",x"58",x"a6",x"cc"),
   752 => (x"66",x"c4",x"7a",x"66"),
   753 => (x"f8",x"49",x"73",x"1e"),
   754 => (x"86",x"c4",x"87",x"f5"),
   755 => (x"1e",x"c8",x"e4",x"c2"),
   756 => (x"f9",x"f9",x"49",x"73"),
   757 => (x"49",x"a3",x"d0",x"87"),
   758 => (x"79",x"66",x"f4",x"c0"),
   759 => (x"26",x"8e",x"dc",x"ff"),
   760 => (x"26",x"4c",x"26",x"4d"),
   761 => (x"0e",x"4f",x"26",x"4b"),
   762 => (x"0e",x"5c",x"5b",x"5e"),
   763 => (x"4b",x"c0",x"4a",x"71"),
   764 => (x"c0",x"02",x"9a",x"72"),
   765 => (x"a2",x"da",x"87",x"e0"),
   766 => (x"4b",x"69",x"9f",x"49"),
   767 => (x"bf",x"d0",x"ec",x"c2"),
   768 => (x"d4",x"87",x"cf",x"02"),
   769 => (x"69",x"9f",x"49",x"a2"),
   770 => (x"ff",x"c0",x"4c",x"49"),
   771 => (x"34",x"d0",x"9c",x"ff"),
   772 => (x"4c",x"c0",x"87",x"c2"),
   773 => (x"9b",x"73",x"b3",x"74"),
   774 => (x"4a",x"87",x"df",x"02"),
   775 => (x"ec",x"c2",x"8a",x"c2"),
   776 => (x"92",x"49",x"bf",x"c8"),
   777 => (x"bf",x"ec",x"f0",x"c2"),
   778 => (x"c2",x"80",x"72",x"48"),
   779 => (x"71",x"58",x"cc",x"f1"),
   780 => (x"c2",x"30",x"c4",x"48"),
   781 => (x"c0",x"58",x"d8",x"ec"),
   782 => (x"f0",x"c2",x"87",x"e9"),
   783 => (x"c2",x"4b",x"bf",x"f0"),
   784 => (x"c2",x"48",x"c8",x"f1"),
   785 => (x"78",x"bf",x"f4",x"f0"),
   786 => (x"bf",x"d0",x"ec",x"c2"),
   787 => (x"c2",x"87",x"c9",x"02"),
   788 => (x"49",x"bf",x"c8",x"ec"),
   789 => (x"87",x"c7",x"31",x"c4"),
   790 => (x"bf",x"f8",x"f0",x"c2"),
   791 => (x"c2",x"31",x"c4",x"49"),
   792 => (x"c2",x"59",x"d8",x"ec"),
   793 => (x"26",x"5b",x"c8",x"f1"),
   794 => (x"26",x"4b",x"26",x"4c"),
   795 => (x"5b",x"5e",x"0e",x"4f"),
   796 => (x"f0",x"0e",x"5d",x"5c"),
   797 => (x"59",x"a6",x"c8",x"86"),
   798 => (x"ff",x"ff",x"ff",x"cf"),
   799 => (x"7e",x"c0",x"4c",x"f8"),
   800 => (x"d8",x"02",x"66",x"c4"),
   801 => (x"c4",x"e4",x"c2",x"87"),
   802 => (x"c2",x"78",x"c0",x"48"),
   803 => (x"c2",x"48",x"fc",x"e3"),
   804 => (x"78",x"bf",x"c8",x"f1"),
   805 => (x"48",x"c0",x"e4",x"c2"),
   806 => (x"bf",x"c4",x"f1",x"c2"),
   807 => (x"e5",x"ec",x"c2",x"78"),
   808 => (x"c2",x"50",x"c0",x"48"),
   809 => (x"49",x"bf",x"d4",x"ec"),
   810 => (x"bf",x"c4",x"e4",x"c2"),
   811 => (x"03",x"aa",x"71",x"4a"),
   812 => (x"72",x"87",x"cc",x"c4"),
   813 => (x"05",x"99",x"cf",x"49"),
   814 => (x"c0",x"87",x"ea",x"c0"),
   815 => (x"c2",x"48",x"e8",x"f9"),
   816 => (x"78",x"bf",x"fc",x"e3"),
   817 => (x"1e",x"c8",x"e4",x"c2"),
   818 => (x"bf",x"fc",x"e3",x"c2"),
   819 => (x"fc",x"e3",x"c2",x"49"),
   820 => (x"78",x"a1",x"c1",x"48"),
   821 => (x"fd",x"df",x"ff",x"71"),
   822 => (x"c0",x"86",x"c4",x"87"),
   823 => (x"c2",x"48",x"e4",x"f9"),
   824 => (x"cc",x"78",x"c8",x"e4"),
   825 => (x"e4",x"f9",x"c0",x"87"),
   826 => (x"e0",x"c0",x"48",x"bf"),
   827 => (x"e8",x"f9",x"c0",x"80"),
   828 => (x"c4",x"e4",x"c2",x"58"),
   829 => (x"80",x"c1",x"48",x"bf"),
   830 => (x"58",x"c8",x"e4",x"c2"),
   831 => (x"00",x"0e",x"64",x"27"),
   832 => (x"bf",x"97",x"bf",x"00"),
   833 => (x"c2",x"02",x"9d",x"4d"),
   834 => (x"e5",x"c3",x"87",x"e5"),
   835 => (x"de",x"c2",x"02",x"ad"),
   836 => (x"e4",x"f9",x"c0",x"87"),
   837 => (x"a3",x"cb",x"4b",x"bf"),
   838 => (x"cf",x"4c",x"11",x"49"),
   839 => (x"d2",x"c1",x"05",x"ac"),
   840 => (x"df",x"49",x"75",x"87"),
   841 => (x"cd",x"89",x"c1",x"99"),
   842 => (x"d8",x"ec",x"c2",x"91"),
   843 => (x"4a",x"a3",x"c1",x"81"),
   844 => (x"a3",x"c3",x"51",x"12"),
   845 => (x"c5",x"51",x"12",x"4a"),
   846 => (x"51",x"12",x"4a",x"a3"),
   847 => (x"12",x"4a",x"a3",x"c7"),
   848 => (x"4a",x"a3",x"c9",x"51"),
   849 => (x"a3",x"ce",x"51",x"12"),
   850 => (x"d0",x"51",x"12",x"4a"),
   851 => (x"51",x"12",x"4a",x"a3"),
   852 => (x"12",x"4a",x"a3",x"d2"),
   853 => (x"4a",x"a3",x"d4",x"51"),
   854 => (x"a3",x"d6",x"51",x"12"),
   855 => (x"d8",x"51",x"12",x"4a"),
   856 => (x"51",x"12",x"4a",x"a3"),
   857 => (x"12",x"4a",x"a3",x"dc"),
   858 => (x"4a",x"a3",x"de",x"51"),
   859 => (x"7e",x"c1",x"51",x"12"),
   860 => (x"74",x"87",x"fc",x"c0"),
   861 => (x"05",x"99",x"c8",x"49"),
   862 => (x"74",x"87",x"ed",x"c0"),
   863 => (x"05",x"99",x"d0",x"49"),
   864 => (x"e0",x"c0",x"87",x"d3"),
   865 => (x"cc",x"c0",x"02",x"66"),
   866 => (x"c0",x"49",x"73",x"87"),
   867 => (x"70",x"0f",x"66",x"e0"),
   868 => (x"d3",x"c0",x"02",x"98"),
   869 => (x"c0",x"05",x"6e",x"87"),
   870 => (x"ec",x"c2",x"87",x"c6"),
   871 => (x"50",x"c0",x"48",x"d8"),
   872 => (x"bf",x"e4",x"f9",x"c0"),
   873 => (x"87",x"eb",x"c2",x"48"),
   874 => (x"48",x"e5",x"ec",x"c2"),
   875 => (x"c2",x"7e",x"50",x"c0"),
   876 => (x"49",x"bf",x"d4",x"ec"),
   877 => (x"bf",x"c4",x"e4",x"c2"),
   878 => (x"04",x"aa",x"71",x"4a"),
   879 => (x"cf",x"87",x"f4",x"fb"),
   880 => (x"f8",x"ff",x"ff",x"ff"),
   881 => (x"c8",x"f1",x"c2",x"4c"),
   882 => (x"c8",x"c0",x"05",x"bf"),
   883 => (x"d0",x"ec",x"c2",x"87"),
   884 => (x"fc",x"c1",x"02",x"bf"),
   885 => (x"c0",x"e4",x"c2",x"87"),
   886 => (x"c4",x"eb",x"49",x"bf"),
   887 => (x"c4",x"e4",x"c2",x"87"),
   888 => (x"48",x"a6",x"c4",x"58"),
   889 => (x"bf",x"c0",x"e4",x"c2"),
   890 => (x"d0",x"ec",x"c2",x"78"),
   891 => (x"db",x"c0",x"02",x"bf"),
   892 => (x"49",x"66",x"c4",x"87"),
   893 => (x"a9",x"74",x"99",x"74"),
   894 => (x"87",x"c8",x"c0",x"02"),
   895 => (x"c0",x"48",x"a6",x"c8"),
   896 => (x"87",x"e7",x"c0",x"78"),
   897 => (x"c1",x"48",x"a6",x"c8"),
   898 => (x"87",x"df",x"c0",x"78"),
   899 => (x"cf",x"49",x"66",x"c4"),
   900 => (x"a9",x"99",x"f8",x"ff"),
   901 => (x"87",x"c8",x"c0",x"02"),
   902 => (x"c0",x"48",x"a6",x"cc"),
   903 => (x"87",x"c5",x"c0",x"78"),
   904 => (x"c1",x"48",x"a6",x"cc"),
   905 => (x"48",x"a6",x"c8",x"78"),
   906 => (x"c8",x"78",x"66",x"cc"),
   907 => (x"e0",x"c0",x"05",x"66"),
   908 => (x"49",x"66",x"c4",x"87"),
   909 => (x"ec",x"c2",x"89",x"c2"),
   910 => (x"91",x"4a",x"bf",x"c8"),
   911 => (x"bf",x"ec",x"f0",x"c2"),
   912 => (x"fc",x"e3",x"c2",x"4a"),
   913 => (x"78",x"a1",x"72",x"48"),
   914 => (x"48",x"c4",x"e4",x"c2"),
   915 => (x"d2",x"f9",x"78",x"c0"),
   916 => (x"cf",x"48",x"c0",x"87"),
   917 => (x"f8",x"ff",x"ff",x"ff"),
   918 => (x"26",x"8e",x"f0",x"4c"),
   919 => (x"26",x"4c",x"26",x"4d"),
   920 => (x"00",x"4f",x"26",x"4b"),
   921 => (x"00",x"00",x"00",x"00"),
   922 => (x"ff",x"ff",x"ff",x"ff"),
   923 => (x"48",x"d4",x"ff",x"1e"),
   924 => (x"68",x"78",x"ff",x"c3"),
   925 => (x"1e",x"4f",x"26",x"48"),
   926 => (x"c3",x"48",x"d4",x"ff"),
   927 => (x"d0",x"ff",x"78",x"ff"),
   928 => (x"78",x"e1",x"c0",x"48"),
   929 => (x"d4",x"48",x"d4",x"ff"),
   930 => (x"1e",x"4f",x"26",x"78"),
   931 => (x"c0",x"48",x"d0",x"ff"),
   932 => (x"4f",x"26",x"78",x"e0"),
   933 => (x"87",x"d4",x"ff",x"1e"),
   934 => (x"02",x"99",x"49",x"70"),
   935 => (x"fb",x"c0",x"87",x"c6"),
   936 => (x"87",x"f1",x"05",x"a9"),
   937 => (x"4f",x"26",x"48",x"71"),
   938 => (x"5c",x"5b",x"5e",x"0e"),
   939 => (x"c0",x"4b",x"71",x"0e"),
   940 => (x"87",x"f8",x"fe",x"4c"),
   941 => (x"02",x"99",x"49",x"70"),
   942 => (x"c0",x"87",x"f9",x"c0"),
   943 => (x"c0",x"02",x"a9",x"ec"),
   944 => (x"fb",x"c0",x"87",x"f2"),
   945 => (x"eb",x"c0",x"02",x"a9"),
   946 => (x"b7",x"66",x"cc",x"87"),
   947 => (x"87",x"c7",x"03",x"ac"),
   948 => (x"c2",x"02",x"66",x"d0"),
   949 => (x"71",x"53",x"71",x"87"),
   950 => (x"87",x"c2",x"02",x"99"),
   951 => (x"cb",x"fe",x"84",x"c1"),
   952 => (x"99",x"49",x"70",x"87"),
   953 => (x"c0",x"87",x"cd",x"02"),
   954 => (x"c7",x"02",x"a9",x"ec"),
   955 => (x"a9",x"fb",x"c0",x"87"),
   956 => (x"87",x"d5",x"ff",x"05"),
   957 => (x"c3",x"02",x"66",x"d0"),
   958 => (x"7b",x"97",x"c0",x"87"),
   959 => (x"05",x"a9",x"fb",x"c0"),
   960 => (x"4a",x"74",x"87",x"c7"),
   961 => (x"c2",x"8a",x"0a",x"c0"),
   962 => (x"72",x"4a",x"74",x"87"),
   963 => (x"26",x"4c",x"26",x"48"),
   964 => (x"1e",x"4f",x"26",x"4b"),
   965 => (x"70",x"87",x"d5",x"fd"),
   966 => (x"f0",x"c0",x"4a",x"49"),
   967 => (x"87",x"c9",x"04",x"aa"),
   968 => (x"01",x"aa",x"f9",x"c0"),
   969 => (x"f0",x"c0",x"87",x"c3"),
   970 => (x"aa",x"c1",x"c1",x"8a"),
   971 => (x"c1",x"87",x"c9",x"04"),
   972 => (x"c3",x"01",x"aa",x"da"),
   973 => (x"8a",x"f7",x"c0",x"87"),
   974 => (x"4f",x"26",x"48",x"72"),
   975 => (x"5c",x"5b",x"5e",x"0e"),
   976 => (x"86",x"f8",x"0e",x"5d"),
   977 => (x"7e",x"c0",x"4c",x"71"),
   978 => (x"c0",x"87",x"ec",x"fc"),
   979 => (x"dc",x"ff",x"c0",x"4b"),
   980 => (x"c0",x"49",x"bf",x"97"),
   981 => (x"87",x"cf",x"04",x"a9"),
   982 => (x"c1",x"87",x"f9",x"fc"),
   983 => (x"dc",x"ff",x"c0",x"83"),
   984 => (x"ab",x"49",x"bf",x"97"),
   985 => (x"c0",x"87",x"f1",x"06"),
   986 => (x"bf",x"97",x"dc",x"ff"),
   987 => (x"fb",x"87",x"cf",x"02"),
   988 => (x"49",x"70",x"87",x"fa"),
   989 => (x"87",x"c6",x"02",x"99"),
   990 => (x"05",x"a9",x"ec",x"c0"),
   991 => (x"4b",x"c0",x"87",x"f1"),
   992 => (x"70",x"87",x"e9",x"fb"),
   993 => (x"87",x"e4",x"fb",x"4d"),
   994 => (x"fb",x"58",x"a6",x"c8"),
   995 => (x"4a",x"70",x"87",x"de"),
   996 => (x"a4",x"c8",x"83",x"c1"),
   997 => (x"49",x"69",x"97",x"49"),
   998 => (x"87",x"da",x"05",x"ad"),
   999 => (x"97",x"49",x"a4",x"c9"),
  1000 => (x"66",x"c4",x"49",x"69"),
  1001 => (x"87",x"ce",x"05",x"a9"),
  1002 => (x"97",x"49",x"a4",x"ca"),
  1003 => (x"05",x"aa",x"49",x"69"),
  1004 => (x"7e",x"c1",x"87",x"c4"),
  1005 => (x"ec",x"c0",x"87",x"d0"),
  1006 => (x"87",x"c6",x"02",x"ad"),
  1007 => (x"05",x"ad",x"fb",x"c0"),
  1008 => (x"4b",x"c0",x"87",x"c4"),
  1009 => (x"02",x"6e",x"7e",x"c1"),
  1010 => (x"fa",x"87",x"f5",x"fe"),
  1011 => (x"48",x"73",x"87",x"fd"),
  1012 => (x"4d",x"26",x"8e",x"f8"),
  1013 => (x"4b",x"26",x"4c",x"26"),
  1014 => (x"00",x"00",x"4f",x"26"),
  1015 => (x"1e",x"73",x"1e",x"00"),
  1016 => (x"c8",x"4b",x"d4",x"ff"),
  1017 => (x"d0",x"ff",x"4a",x"66"),
  1018 => (x"78",x"c5",x"c8",x"48"),
  1019 => (x"c1",x"48",x"d4",x"ff"),
  1020 => (x"7b",x"11",x"78",x"d4"),
  1021 => (x"f9",x"05",x"8a",x"c1"),
  1022 => (x"48",x"d0",x"ff",x"87"),
  1023 => (x"4b",x"26",x"78",x"c4"),
  1024 => (x"5e",x"0e",x"4f",x"26"),
  1025 => (x"0e",x"5d",x"5c",x"5b"),
  1026 => (x"7e",x"71",x"86",x"f8"),
  1027 => (x"f1",x"c2",x"1e",x"6e"),
  1028 => (x"c3",x"e4",x"49",x"dc"),
  1029 => (x"70",x"86",x"c4",x"87"),
  1030 => (x"e4",x"c4",x"02",x"98"),
  1031 => (x"f4",x"ec",x"c1",x"87"),
  1032 => (x"49",x"6e",x"4c",x"bf"),
  1033 => (x"c8",x"87",x"d5",x"fc"),
  1034 => (x"98",x"70",x"58",x"a6"),
  1035 => (x"c4",x"87",x"c5",x"05"),
  1036 => (x"78",x"c1",x"48",x"a6"),
  1037 => (x"c5",x"48",x"d0",x"ff"),
  1038 => (x"48",x"d4",x"ff",x"78"),
  1039 => (x"c4",x"78",x"d5",x"c1"),
  1040 => (x"89",x"c1",x"49",x"66"),
  1041 => (x"ec",x"c1",x"31",x"c6"),
  1042 => (x"4a",x"bf",x"97",x"ec"),
  1043 => (x"ff",x"b0",x"71",x"48"),
  1044 => (x"ff",x"78",x"08",x"d4"),
  1045 => (x"78",x"c4",x"48",x"d0"),
  1046 => (x"97",x"d8",x"f1",x"c2"),
  1047 => (x"99",x"d0",x"49",x"bf"),
  1048 => (x"c5",x"87",x"dd",x"02"),
  1049 => (x"48",x"d4",x"ff",x"78"),
  1050 => (x"c0",x"78",x"d6",x"c1"),
  1051 => (x"48",x"d4",x"ff",x"4a"),
  1052 => (x"c1",x"78",x"ff",x"c3"),
  1053 => (x"aa",x"e0",x"c0",x"82"),
  1054 => (x"ff",x"87",x"f2",x"04"),
  1055 => (x"78",x"c4",x"48",x"d0"),
  1056 => (x"c3",x"48",x"d4",x"ff"),
  1057 => (x"d0",x"ff",x"78",x"ff"),
  1058 => (x"ff",x"78",x"c5",x"48"),
  1059 => (x"d3",x"c1",x"48",x"d4"),
  1060 => (x"ff",x"78",x"c1",x"78"),
  1061 => (x"78",x"c4",x"48",x"d0"),
  1062 => (x"06",x"ac",x"b7",x"c0"),
  1063 => (x"c2",x"87",x"cb",x"c2"),
  1064 => (x"4b",x"bf",x"e4",x"f1"),
  1065 => (x"73",x"7e",x"74",x"8c"),
  1066 => (x"dd",x"c1",x"02",x"9b"),
  1067 => (x"4d",x"c0",x"c8",x"87"),
  1068 => (x"ab",x"b7",x"c0",x"8b"),
  1069 => (x"c8",x"87",x"c6",x"03"),
  1070 => (x"c0",x"4d",x"a3",x"c0"),
  1071 => (x"d8",x"f1",x"c2",x"4b"),
  1072 => (x"d0",x"49",x"bf",x"97"),
  1073 => (x"87",x"cf",x"02",x"99"),
  1074 => (x"f1",x"c2",x"1e",x"c0"),
  1075 => (x"fd",x"e5",x"49",x"dc"),
  1076 => (x"70",x"86",x"c4",x"87"),
  1077 => (x"c2",x"87",x"d8",x"4c"),
  1078 => (x"c2",x"1e",x"c8",x"e4"),
  1079 => (x"e5",x"49",x"dc",x"f1"),
  1080 => (x"4c",x"70",x"87",x"ec"),
  1081 => (x"e4",x"c2",x"1e",x"75"),
  1082 => (x"f0",x"fb",x"49",x"c8"),
  1083 => (x"74",x"86",x"c8",x"87"),
  1084 => (x"87",x"c5",x"05",x"9c"),
  1085 => (x"ca",x"c1",x"48",x"c0"),
  1086 => (x"c2",x"1e",x"c1",x"87"),
  1087 => (x"e3",x"49",x"dc",x"f1"),
  1088 => (x"86",x"c4",x"87",x"fd"),
  1089 => (x"fe",x"05",x"9b",x"73"),
  1090 => (x"4c",x"6e",x"87",x"e3"),
  1091 => (x"06",x"ac",x"b7",x"c0"),
  1092 => (x"f1",x"c2",x"87",x"d1"),
  1093 => (x"78",x"c0",x"48",x"dc"),
  1094 => (x"78",x"c0",x"80",x"d0"),
  1095 => (x"f1",x"c2",x"80",x"f4"),
  1096 => (x"c0",x"78",x"bf",x"e8"),
  1097 => (x"fd",x"01",x"ac",x"b7"),
  1098 => (x"d0",x"ff",x"87",x"f5"),
  1099 => (x"ff",x"78",x"c5",x"48"),
  1100 => (x"d3",x"c1",x"48",x"d4"),
  1101 => (x"ff",x"78",x"c0",x"78"),
  1102 => (x"78",x"c4",x"48",x"d0"),
  1103 => (x"c2",x"c0",x"48",x"c1"),
  1104 => (x"f8",x"48",x"c0",x"87"),
  1105 => (x"26",x"4d",x"26",x"8e"),
  1106 => (x"26",x"4b",x"26",x"4c"),
  1107 => (x"5b",x"5e",x"0e",x"4f"),
  1108 => (x"fc",x"0e",x"5d",x"5c"),
  1109 => (x"c0",x"4d",x"71",x"86"),
  1110 => (x"04",x"ad",x"4c",x"4b"),
  1111 => (x"c0",x"87",x"e8",x"c0"),
  1112 => (x"74",x"1e",x"fc",x"fc"),
  1113 => (x"87",x"c4",x"02",x"9c"),
  1114 => (x"87",x"c2",x"4a",x"c0"),
  1115 => (x"49",x"72",x"4a",x"c1"),
  1116 => (x"c4",x"87",x"fa",x"eb"),
  1117 => (x"c1",x"7e",x"70",x"86"),
  1118 => (x"c2",x"05",x"6e",x"83"),
  1119 => (x"c1",x"4b",x"75",x"87"),
  1120 => (x"06",x"ab",x"75",x"84"),
  1121 => (x"6e",x"87",x"d8",x"ff"),
  1122 => (x"26",x"8e",x"fc",x"48"),
  1123 => (x"26",x"4c",x"26",x"4d"),
  1124 => (x"0e",x"4f",x"26",x"4b"),
  1125 => (x"0e",x"5c",x"5b",x"5e"),
  1126 => (x"66",x"cc",x"4b",x"71"),
  1127 => (x"4c",x"87",x"d8",x"02"),
  1128 => (x"02",x"8c",x"f0",x"c0"),
  1129 => (x"4a",x"74",x"87",x"d8"),
  1130 => (x"d1",x"02",x"8a",x"c1"),
  1131 => (x"cd",x"02",x"8a",x"87"),
  1132 => (x"c9",x"02",x"8a",x"87"),
  1133 => (x"73",x"87",x"d9",x"87"),
  1134 => (x"87",x"c6",x"f9",x"49"),
  1135 => (x"1e",x"74",x"87",x"d2"),
  1136 => (x"d9",x"c1",x"49",x"c0"),
  1137 => (x"1e",x"74",x"87",x"ca"),
  1138 => (x"d9",x"c1",x"49",x"73"),
  1139 => (x"86",x"c8",x"87",x"c2"),
  1140 => (x"4b",x"26",x"4c",x"26"),
  1141 => (x"5e",x"0e",x"4f",x"26"),
  1142 => (x"0e",x"5d",x"5c",x"5b"),
  1143 => (x"4c",x"71",x"86",x"fc"),
  1144 => (x"c2",x"91",x"de",x"49"),
  1145 => (x"71",x"4d",x"fc",x"f2"),
  1146 => (x"02",x"6d",x"97",x"85"),
  1147 => (x"c2",x"87",x"dc",x"c1"),
  1148 => (x"49",x"bf",x"ec",x"f2"),
  1149 => (x"fd",x"71",x"81",x"74"),
  1150 => (x"7e",x"70",x"87",x"d3"),
  1151 => (x"c0",x"02",x"98",x"48"),
  1152 => (x"f2",x"c2",x"87",x"f2"),
  1153 => (x"4a",x"70",x"4b",x"f0"),
  1154 => (x"fb",x"fe",x"49",x"cb"),
  1155 => (x"4b",x"74",x"87",x"f2"),
  1156 => (x"ec",x"c1",x"93",x"cc"),
  1157 => (x"83",x"c4",x"83",x"f8"),
  1158 => (x"7b",x"d8",x"c9",x"c1"),
  1159 => (x"c2",x"c1",x"49",x"74"),
  1160 => (x"7b",x"75",x"87",x"ea"),
  1161 => (x"97",x"f0",x"ec",x"c1"),
  1162 => (x"c2",x"1e",x"49",x"bf"),
  1163 => (x"fd",x"49",x"f0",x"f2"),
  1164 => (x"86",x"c4",x"87",x"e1"),
  1165 => (x"c2",x"c1",x"49",x"74"),
  1166 => (x"49",x"c0",x"87",x"d2"),
  1167 => (x"87",x"ed",x"c3",x"c1"),
  1168 => (x"48",x"d4",x"f1",x"c2"),
  1169 => (x"c0",x"49",x"50",x"c0"),
  1170 => (x"fc",x"87",x"c5",x"e1"),
  1171 => (x"26",x"4d",x"26",x"8e"),
  1172 => (x"26",x"4b",x"26",x"4c"),
  1173 => (x"00",x"00",x"00",x"4f"),
  1174 => (x"64",x"61",x"6f",x"4c"),
  1175 => (x"2e",x"67",x"6e",x"69"),
  1176 => (x"00",x"00",x"2e",x"2e"),
  1177 => (x"61",x"42",x"20",x"80"),
  1178 => (x"00",x"00",x"6b",x"63"),
  1179 => (x"64",x"61",x"6f",x"4c"),
  1180 => (x"20",x"2e",x"2a",x"20"),
  1181 => (x"00",x"00",x"00",x"00"),
  1182 => (x"00",x"00",x"20",x"3a"),
  1183 => (x"61",x"42",x"20",x"80"),
  1184 => (x"00",x"00",x"6b",x"63"),
  1185 => (x"78",x"45",x"20",x"80"),
  1186 => (x"00",x"00",x"74",x"69"),
  1187 => (x"49",x"20",x"44",x"53"),
  1188 => (x"2e",x"74",x"69",x"6e"),
  1189 => (x"00",x"00",x"00",x"2e"),
  1190 => (x"00",x"00",x"4b",x"4f"),
  1191 => (x"54",x"4f",x"4f",x"42"),
  1192 => (x"20",x"20",x"20",x"20"),
  1193 => (x"00",x"4d",x"4f",x"52"),
  1194 => (x"71",x"1e",x"73",x"1e"),
  1195 => (x"f2",x"c2",x"49",x"4b"),
  1196 => (x"71",x"81",x"bf",x"ec"),
  1197 => (x"70",x"87",x"d6",x"fa"),
  1198 => (x"c4",x"02",x"9a",x"4a"),
  1199 => (x"e6",x"e4",x"49",x"87"),
  1200 => (x"ec",x"f2",x"c2",x"87"),
  1201 => (x"73",x"78",x"c0",x"48"),
  1202 => (x"87",x"fa",x"c1",x"49"),
  1203 => (x"4f",x"26",x"4b",x"26"),
  1204 => (x"71",x"1e",x"73",x"1e"),
  1205 => (x"4a",x"a3",x"c4",x"4b"),
  1206 => (x"87",x"d0",x"c1",x"02"),
  1207 => (x"dc",x"02",x"8a",x"c1"),
  1208 => (x"c0",x"02",x"8a",x"87"),
  1209 => (x"05",x"8a",x"87",x"f2"),
  1210 => (x"c2",x"87",x"d3",x"c1"),
  1211 => (x"02",x"bf",x"ec",x"f2"),
  1212 => (x"48",x"87",x"cb",x"c1"),
  1213 => (x"f2",x"c2",x"88",x"c1"),
  1214 => (x"c1",x"c1",x"58",x"f0"),
  1215 => (x"ec",x"f2",x"c2",x"87"),
  1216 => (x"89",x"c6",x"49",x"bf"),
  1217 => (x"59",x"f0",x"f2",x"c2"),
  1218 => (x"03",x"a9",x"b7",x"c0"),
  1219 => (x"c2",x"87",x"ef",x"c0"),
  1220 => (x"c0",x"48",x"ec",x"f2"),
  1221 => (x"87",x"e6",x"c0",x"78"),
  1222 => (x"bf",x"e8",x"f2",x"c2"),
  1223 => (x"c2",x"87",x"df",x"02"),
  1224 => (x"48",x"bf",x"ec",x"f2"),
  1225 => (x"f2",x"c2",x"80",x"c1"),
  1226 => (x"87",x"d2",x"58",x"f0"),
  1227 => (x"bf",x"e8",x"f2",x"c2"),
  1228 => (x"c2",x"87",x"cb",x"02"),
  1229 => (x"48",x"bf",x"ec",x"f2"),
  1230 => (x"f2",x"c2",x"80",x"c6"),
  1231 => (x"49",x"73",x"58",x"f0"),
  1232 => (x"4b",x"26",x"87",x"c4"),
  1233 => (x"5e",x"0e",x"4f",x"26"),
  1234 => (x"0e",x"5d",x"5c",x"5b"),
  1235 => (x"a6",x"d0",x"86",x"f0"),
  1236 => (x"c8",x"e4",x"c2",x"59"),
  1237 => (x"c2",x"4c",x"c0",x"4d"),
  1238 => (x"c1",x"48",x"e8",x"f2"),
  1239 => (x"48",x"a6",x"c4",x"78"),
  1240 => (x"7e",x"75",x"78",x"c0"),
  1241 => (x"bf",x"ec",x"f2",x"c2"),
  1242 => (x"06",x"a8",x"c0",x"48"),
  1243 => (x"75",x"87",x"fa",x"c0"),
  1244 => (x"c8",x"e4",x"c2",x"7e"),
  1245 => (x"c0",x"02",x"98",x"48"),
  1246 => (x"fc",x"c0",x"87",x"ef"),
  1247 => (x"66",x"c8",x"1e",x"fc"),
  1248 => (x"c0",x"87",x"c4",x"02"),
  1249 => (x"c1",x"87",x"c2",x"4d"),
  1250 => (x"e3",x"49",x"75",x"4d"),
  1251 => (x"86",x"c4",x"87",x"df"),
  1252 => (x"84",x"c1",x"7e",x"70"),
  1253 => (x"c1",x"48",x"66",x"c4"),
  1254 => (x"58",x"a6",x"c8",x"80"),
  1255 => (x"bf",x"ec",x"f2",x"c2"),
  1256 => (x"87",x"c5",x"03",x"ac"),
  1257 => (x"d1",x"ff",x"05",x"6e"),
  1258 => (x"c0",x"4d",x"6e",x"87"),
  1259 => (x"02",x"9d",x"75",x"4c"),
  1260 => (x"c0",x"87",x"e0",x"c3"),
  1261 => (x"c8",x"1e",x"fc",x"fc"),
  1262 => (x"87",x"c7",x"02",x"66"),
  1263 => (x"c0",x"48",x"a6",x"cc"),
  1264 => (x"cc",x"87",x"c5",x"78"),
  1265 => (x"78",x"c1",x"48",x"a6"),
  1266 => (x"e2",x"49",x"66",x"cc"),
  1267 => (x"86",x"c4",x"87",x"df"),
  1268 => (x"98",x"48",x"7e",x"70"),
  1269 => (x"87",x"e8",x"c2",x"02"),
  1270 => (x"97",x"81",x"cb",x"49"),
  1271 => (x"99",x"d0",x"49",x"69"),
  1272 => (x"87",x"d6",x"c1",x"02"),
  1273 => (x"4a",x"e8",x"ca",x"c1"),
  1274 => (x"91",x"cc",x"49",x"74"),
  1275 => (x"81",x"f8",x"ec",x"c1"),
  1276 => (x"81",x"c8",x"79",x"72"),
  1277 => (x"74",x"51",x"ff",x"c3"),
  1278 => (x"c2",x"91",x"de",x"49"),
  1279 => (x"71",x"4d",x"fc",x"f2"),
  1280 => (x"97",x"c1",x"c2",x"85"),
  1281 => (x"49",x"a5",x"c1",x"7d"),
  1282 => (x"c2",x"51",x"e0",x"c0"),
  1283 => (x"bf",x"97",x"d8",x"ec"),
  1284 => (x"c1",x"87",x"d2",x"02"),
  1285 => (x"4b",x"a5",x"c2",x"84"),
  1286 => (x"4a",x"d8",x"ec",x"c2"),
  1287 => (x"f3",x"fe",x"49",x"db"),
  1288 => (x"db",x"c1",x"87",x"de"),
  1289 => (x"49",x"a5",x"cd",x"87"),
  1290 => (x"84",x"c1",x"51",x"c0"),
  1291 => (x"6e",x"4b",x"a5",x"c2"),
  1292 => (x"fe",x"49",x"cb",x"4a"),
  1293 => (x"c1",x"87",x"c9",x"f3"),
  1294 => (x"c7",x"c1",x"87",x"c6"),
  1295 => (x"49",x"74",x"4a",x"d6"),
  1296 => (x"ec",x"c1",x"91",x"cc"),
  1297 => (x"79",x"72",x"81",x"f8"),
  1298 => (x"97",x"d8",x"ec",x"c2"),
  1299 => (x"87",x"d8",x"02",x"bf"),
  1300 => (x"91",x"de",x"49",x"74"),
  1301 => (x"f2",x"c2",x"84",x"c1"),
  1302 => (x"83",x"71",x"4b",x"fc"),
  1303 => (x"4a",x"d8",x"ec",x"c2"),
  1304 => (x"f2",x"fe",x"49",x"dd"),
  1305 => (x"87",x"d8",x"87",x"da"),
  1306 => (x"93",x"de",x"4b",x"74"),
  1307 => (x"83",x"fc",x"f2",x"c2"),
  1308 => (x"c0",x"49",x"a3",x"cb"),
  1309 => (x"73",x"84",x"c1",x"51"),
  1310 => (x"49",x"cb",x"4a",x"6e"),
  1311 => (x"87",x"c0",x"f2",x"fe"),
  1312 => (x"c1",x"48",x"66",x"c4"),
  1313 => (x"58",x"a6",x"c8",x"80"),
  1314 => (x"c0",x"03",x"ac",x"c7"),
  1315 => (x"05",x"6e",x"87",x"c5"),
  1316 => (x"c7",x"87",x"e0",x"fc"),
  1317 => (x"e6",x"c0",x"03",x"ac"),
  1318 => (x"e8",x"f2",x"c2",x"87"),
  1319 => (x"c1",x"78",x"c0",x"48"),
  1320 => (x"74",x"4a",x"d6",x"c7"),
  1321 => (x"c1",x"91",x"cc",x"49"),
  1322 => (x"72",x"81",x"f8",x"ec"),
  1323 => (x"de",x"49",x"74",x"79"),
  1324 => (x"fc",x"f2",x"c2",x"91"),
  1325 => (x"c1",x"51",x"c0",x"81"),
  1326 => (x"04",x"ac",x"c7",x"84"),
  1327 => (x"c1",x"87",x"da",x"ff"),
  1328 => (x"c0",x"48",x"d4",x"ee"),
  1329 => (x"c1",x"80",x"f7",x"50"),
  1330 => (x"c1",x"40",x"ec",x"d4"),
  1331 => (x"c8",x"78",x"e4",x"c9"),
  1332 => (x"d0",x"cb",x"c1",x"80"),
  1333 => (x"49",x"66",x"cc",x"78"),
  1334 => (x"87",x"f0",x"f7",x"c0"),
  1335 => (x"4d",x"26",x"8e",x"f0"),
  1336 => (x"4b",x"26",x"4c",x"26"),
  1337 => (x"73",x"1e",x"4f",x"26"),
  1338 => (x"49",x"4b",x"71",x"1e"),
  1339 => (x"ec",x"c1",x"91",x"cc"),
  1340 => (x"a1",x"c8",x"81",x"f8"),
  1341 => (x"ec",x"ec",x"c1",x"4a"),
  1342 => (x"c9",x"50",x"12",x"48"),
  1343 => (x"ff",x"c0",x"4a",x"a1"),
  1344 => (x"50",x"12",x"48",x"dc"),
  1345 => (x"ec",x"c1",x"81",x"ca"),
  1346 => (x"50",x"11",x"48",x"f0"),
  1347 => (x"97",x"f0",x"ec",x"c1"),
  1348 => (x"c0",x"1e",x"49",x"bf"),
  1349 => (x"87",x"fb",x"f1",x"49"),
  1350 => (x"e9",x"f8",x"49",x"73"),
  1351 => (x"26",x"8e",x"fc",x"87"),
  1352 => (x"1e",x"4f",x"26",x"4b"),
  1353 => (x"f8",x"c0",x"49",x"c0"),
  1354 => (x"4f",x"26",x"87",x"c3"),
  1355 => (x"49",x"4a",x"71",x"1e"),
  1356 => (x"ec",x"c1",x"91",x"cc"),
  1357 => (x"81",x"c8",x"81",x"f8"),
  1358 => (x"48",x"d4",x"f1",x"c2"),
  1359 => (x"f0",x"c0",x"50",x"11"),
  1360 => (x"ed",x"fe",x"49",x"a2"),
  1361 => (x"49",x"c0",x"87",x"c6"),
  1362 => (x"26",x"87",x"c5",x"d5"),
  1363 => (x"d4",x"ff",x"1e",x"4f"),
  1364 => (x"7a",x"ff",x"c3",x"4a"),
  1365 => (x"c0",x"48",x"d0",x"ff"),
  1366 => (x"7a",x"de",x"78",x"e1"),
  1367 => (x"c8",x"48",x"7a",x"71"),
  1368 => (x"7a",x"70",x"28",x"b7"),
  1369 => (x"b7",x"d0",x"48",x"71"),
  1370 => (x"71",x"7a",x"70",x"28"),
  1371 => (x"28",x"b7",x"d8",x"48"),
  1372 => (x"d0",x"ff",x"7a",x"70"),
  1373 => (x"78",x"e0",x"c0",x"48"),
  1374 => (x"5e",x"0e",x"4f",x"26"),
  1375 => (x"0e",x"5d",x"5c",x"5b"),
  1376 => (x"4d",x"71",x"86",x"f4"),
  1377 => (x"c1",x"91",x"cc",x"49"),
  1378 => (x"c8",x"81",x"f8",x"ec"),
  1379 => (x"a1",x"ca",x"4a",x"a1"),
  1380 => (x"48",x"a6",x"c4",x"7e"),
  1381 => (x"bf",x"d0",x"f1",x"c2"),
  1382 => (x"bf",x"97",x"6e",x"78"),
  1383 => (x"4c",x"66",x"c4",x"4b"),
  1384 => (x"48",x"12",x"2c",x"73"),
  1385 => (x"70",x"58",x"a6",x"cc"),
  1386 => (x"c9",x"84",x"c1",x"9c"),
  1387 => (x"49",x"69",x"97",x"81"),
  1388 => (x"c2",x"04",x"ac",x"b7"),
  1389 => (x"6e",x"4c",x"c0",x"87"),
  1390 => (x"c8",x"4a",x"bf",x"97"),
  1391 => (x"31",x"72",x"49",x"66"),
  1392 => (x"66",x"c4",x"b9",x"ff"),
  1393 => (x"72",x"48",x"74",x"99"),
  1394 => (x"b1",x"4a",x"70",x"30"),
  1395 => (x"59",x"d4",x"f1",x"c2"),
  1396 => (x"87",x"f9",x"fd",x"71"),
  1397 => (x"f2",x"c2",x"1e",x"c7"),
  1398 => (x"c1",x"1e",x"bf",x"e4"),
  1399 => (x"c2",x"1e",x"f8",x"ec"),
  1400 => (x"bf",x"97",x"d4",x"f1"),
  1401 => (x"87",x"f4",x"c1",x"49"),
  1402 => (x"f3",x"c0",x"49",x"75"),
  1403 => (x"8e",x"e8",x"87",x"de"),
  1404 => (x"4c",x"26",x"4d",x"26"),
  1405 => (x"4f",x"26",x"4b",x"26"),
  1406 => (x"71",x"1e",x"73",x"1e"),
  1407 => (x"f9",x"fd",x"49",x"4b"),
  1408 => (x"fd",x"49",x"73",x"87"),
  1409 => (x"4b",x"26",x"87",x"f4"),
  1410 => (x"73",x"1e",x"4f",x"26"),
  1411 => (x"c2",x"4b",x"71",x"1e"),
  1412 => (x"d6",x"02",x"4a",x"a3"),
  1413 => (x"05",x"8a",x"c1",x"87"),
  1414 => (x"c2",x"87",x"e2",x"c0"),
  1415 => (x"02",x"bf",x"e4",x"f2"),
  1416 => (x"c1",x"48",x"87",x"db"),
  1417 => (x"e8",x"f2",x"c2",x"88"),
  1418 => (x"c2",x"87",x"d2",x"58"),
  1419 => (x"02",x"bf",x"e8",x"f2"),
  1420 => (x"f2",x"c2",x"87",x"cb"),
  1421 => (x"c1",x"48",x"bf",x"e4"),
  1422 => (x"e8",x"f2",x"c2",x"80"),
  1423 => (x"c2",x"1e",x"c7",x"58"),
  1424 => (x"1e",x"bf",x"e4",x"f2"),
  1425 => (x"1e",x"f8",x"ec",x"c1"),
  1426 => (x"97",x"d4",x"f1",x"c2"),
  1427 => (x"87",x"cc",x"49",x"bf"),
  1428 => (x"f1",x"c0",x"49",x"73"),
  1429 => (x"8e",x"f4",x"87",x"f6"),
  1430 => (x"4f",x"26",x"4b",x"26"),
  1431 => (x"5c",x"5b",x"5e",x"0e"),
  1432 => (x"cc",x"ff",x"0e",x"5d"),
  1433 => (x"a6",x"e8",x"c0",x"86"),
  1434 => (x"48",x"a6",x"cc",x"59"),
  1435 => (x"80",x"c4",x"78",x"c0"),
  1436 => (x"80",x"c4",x"78",x"c0"),
  1437 => (x"80",x"c4",x"78",x"c0"),
  1438 => (x"78",x"66",x"c8",x"c1"),
  1439 => (x"78",x"c1",x"80",x"c4"),
  1440 => (x"78",x"c1",x"80",x"c4"),
  1441 => (x"48",x"e8",x"f2",x"c2"),
  1442 => (x"df",x"ff",x"78",x"c1"),
  1443 => (x"c3",x"e0",x"87",x"e9"),
  1444 => (x"d7",x"df",x"ff",x"87"),
  1445 => (x"c0",x"4d",x"70",x"87"),
  1446 => (x"c1",x"02",x"ad",x"fb"),
  1447 => (x"e4",x"c0",x"87",x"f3"),
  1448 => (x"e8",x"c1",x"05",x"66"),
  1449 => (x"66",x"c4",x"c1",x"87"),
  1450 => (x"6a",x"82",x"c4",x"4a"),
  1451 => (x"ec",x"c9",x"c1",x"7e"),
  1452 => (x"20",x"49",x"6e",x"48"),
  1453 => (x"10",x"41",x"20",x"41"),
  1454 => (x"66",x"c4",x"c1",x"51"),
  1455 => (x"e6",x"d3",x"c1",x"48"),
  1456 => (x"c7",x"49",x"6a",x"78"),
  1457 => (x"c1",x"51",x"75",x"81"),
  1458 => (x"c8",x"49",x"66",x"c4"),
  1459 => (x"dc",x"51",x"c1",x"81"),
  1460 => (x"78",x"c2",x"48",x"a6"),
  1461 => (x"49",x"66",x"c4",x"c1"),
  1462 => (x"51",x"c0",x"81",x"c9"),
  1463 => (x"49",x"66",x"c4",x"c1"),
  1464 => (x"51",x"c0",x"81",x"ca"),
  1465 => (x"1e",x"d8",x"1e",x"c1"),
  1466 => (x"81",x"c8",x"49",x"6a"),
  1467 => (x"87",x"f8",x"de",x"ff"),
  1468 => (x"c8",x"c1",x"86",x"c8"),
  1469 => (x"a8",x"c0",x"48",x"66"),
  1470 => (x"d4",x"87",x"c7",x"01"),
  1471 => (x"78",x"c1",x"48",x"a6"),
  1472 => (x"c8",x"c1",x"87",x"cf"),
  1473 => (x"88",x"c1",x"48",x"66"),
  1474 => (x"c4",x"58",x"a6",x"dc"),
  1475 => (x"c3",x"de",x"ff",x"87"),
  1476 => (x"02",x"9d",x"75",x"87"),
  1477 => (x"d4",x"87",x"f1",x"cb"),
  1478 => (x"cc",x"c1",x"48",x"66"),
  1479 => (x"cb",x"03",x"a8",x"66"),
  1480 => (x"7e",x"c0",x"87",x"e6"),
  1481 => (x"87",x"c4",x"dd",x"ff"),
  1482 => (x"c1",x"48",x"4d",x"70"),
  1483 => (x"a6",x"c8",x"88",x"c6"),
  1484 => (x"02",x"98",x"70",x"58"),
  1485 => (x"48",x"87",x"d6",x"c1"),
  1486 => (x"a6",x"c8",x"88",x"c9"),
  1487 => (x"02",x"98",x"70",x"58"),
  1488 => (x"48",x"87",x"d7",x"c5"),
  1489 => (x"a6",x"c8",x"88",x"c1"),
  1490 => (x"02",x"98",x"70",x"58"),
  1491 => (x"48",x"87",x"f8",x"c2"),
  1492 => (x"a6",x"c8",x"88",x"c3"),
  1493 => (x"02",x"98",x"70",x"58"),
  1494 => (x"c1",x"48",x"87",x"cf"),
  1495 => (x"58",x"a6",x"c8",x"88"),
  1496 => (x"c4",x"02",x"98",x"70"),
  1497 => (x"fe",x"c9",x"87",x"f4"),
  1498 => (x"7e",x"f0",x"c0",x"87"),
  1499 => (x"87",x"fc",x"db",x"ff"),
  1500 => (x"ec",x"c0",x"4d",x"70"),
  1501 => (x"87",x"c2",x"02",x"ad"),
  1502 => (x"ec",x"c0",x"7e",x"75"),
  1503 => (x"87",x"cd",x"02",x"ad"),
  1504 => (x"87",x"e8",x"db",x"ff"),
  1505 => (x"ec",x"c0",x"4d",x"70"),
  1506 => (x"f3",x"ff",x"05",x"ad"),
  1507 => (x"66",x"e4",x"c0",x"87"),
  1508 => (x"87",x"ea",x"c1",x"05"),
  1509 => (x"02",x"ad",x"ec",x"c0"),
  1510 => (x"db",x"ff",x"87",x"c4"),
  1511 => (x"1e",x"c0",x"87",x"ce"),
  1512 => (x"66",x"dc",x"1e",x"ca"),
  1513 => (x"c1",x"93",x"cc",x"4b"),
  1514 => (x"c4",x"83",x"66",x"cc"),
  1515 => (x"49",x"6c",x"4c",x"a3"),
  1516 => (x"87",x"f4",x"db",x"ff"),
  1517 => (x"1e",x"de",x"1e",x"c1"),
  1518 => (x"db",x"ff",x"49",x"6c"),
  1519 => (x"86",x"d0",x"87",x"ea"),
  1520 => (x"7b",x"e6",x"d3",x"c1"),
  1521 => (x"dc",x"49",x"a3",x"c8"),
  1522 => (x"a3",x"c9",x"51",x"66"),
  1523 => (x"66",x"e0",x"c0",x"49"),
  1524 => (x"49",x"a3",x"ca",x"51"),
  1525 => (x"66",x"dc",x"51",x"6e"),
  1526 => (x"c0",x"80",x"c1",x"48"),
  1527 => (x"d4",x"58",x"a6",x"e0"),
  1528 => (x"66",x"d8",x"48",x"66"),
  1529 => (x"87",x"cb",x"04",x"a8"),
  1530 => (x"c1",x"48",x"66",x"d4"),
  1531 => (x"58",x"a6",x"d8",x"80"),
  1532 => (x"d8",x"87",x"fa",x"c7"),
  1533 => (x"88",x"c1",x"48",x"66"),
  1534 => (x"c7",x"58",x"a6",x"dc"),
  1535 => (x"da",x"ff",x"87",x"ef"),
  1536 => (x"4d",x"70",x"87",x"d2"),
  1537 => (x"ff",x"87",x"e6",x"c7"),
  1538 => (x"d0",x"87",x"c8",x"dc"),
  1539 => (x"66",x"d0",x"58",x"a6"),
  1540 => (x"87",x"c6",x"06",x"a8"),
  1541 => (x"cc",x"48",x"a6",x"d0"),
  1542 => (x"db",x"ff",x"78",x"66"),
  1543 => (x"ec",x"c0",x"87",x"f5"),
  1544 => (x"f5",x"c1",x"05",x"a8"),
  1545 => (x"66",x"e4",x"c0",x"87"),
  1546 => (x"87",x"e5",x"c1",x"05"),
  1547 => (x"cc",x"49",x"66",x"d4"),
  1548 => (x"66",x"c4",x"c1",x"91"),
  1549 => (x"4a",x"a1",x"c4",x"81"),
  1550 => (x"a1",x"c8",x"4c",x"6a"),
  1551 => (x"52",x"66",x"cc",x"4a"),
  1552 => (x"79",x"ec",x"d4",x"c1"),
  1553 => (x"87",x"e4",x"d8",x"ff"),
  1554 => (x"02",x"9d",x"4d",x"70"),
  1555 => (x"fb",x"c0",x"87",x"da"),
  1556 => (x"87",x"d4",x"02",x"ad"),
  1557 => (x"d8",x"ff",x"54",x"75"),
  1558 => (x"4d",x"70",x"87",x"d2"),
  1559 => (x"c7",x"c0",x"02",x"9d"),
  1560 => (x"ad",x"fb",x"c0",x"87"),
  1561 => (x"87",x"ec",x"ff",x"05"),
  1562 => (x"c2",x"54",x"e0",x"c0"),
  1563 => (x"97",x"c0",x"54",x"c1"),
  1564 => (x"48",x"66",x"d4",x"7c"),
  1565 => (x"04",x"a8",x"66",x"d8"),
  1566 => (x"d4",x"87",x"cb",x"c0"),
  1567 => (x"80",x"c1",x"48",x"66"),
  1568 => (x"c5",x"58",x"a6",x"d8"),
  1569 => (x"66",x"d8",x"87",x"e7"),
  1570 => (x"dc",x"88",x"c1",x"48"),
  1571 => (x"dc",x"c5",x"58",x"a6"),
  1572 => (x"ff",x"d7",x"ff",x"87"),
  1573 => (x"c5",x"4d",x"70",x"87"),
  1574 => (x"66",x"cc",x"87",x"d3"),
  1575 => (x"66",x"e4",x"c0",x"48"),
  1576 => (x"f4",x"c4",x"05",x"a8"),
  1577 => (x"a6",x"e8",x"c0",x"87"),
  1578 => (x"ff",x"78",x"c0",x"48"),
  1579 => (x"70",x"87",x"e4",x"d9"),
  1580 => (x"de",x"d9",x"ff",x"7e"),
  1581 => (x"a6",x"f0",x"c0",x"87"),
  1582 => (x"a8",x"ec",x"c0",x"58"),
  1583 => (x"87",x"c7",x"c0",x"05"),
  1584 => (x"78",x"6e",x"48",x"a6"),
  1585 => (x"ff",x"87",x"c4",x"c0"),
  1586 => (x"d4",x"87",x"e1",x"d6"),
  1587 => (x"91",x"cc",x"49",x"66"),
  1588 => (x"48",x"66",x"c4",x"c1"),
  1589 => (x"a6",x"c8",x"80",x"71"),
  1590 => (x"4a",x"66",x"c4",x"58"),
  1591 => (x"66",x"c4",x"82",x"c8"),
  1592 => (x"6e",x"81",x"ca",x"49"),
  1593 => (x"66",x"ec",x"c0",x"51"),
  1594 => (x"6e",x"81",x"c1",x"49"),
  1595 => (x"71",x"48",x"c1",x"89"),
  1596 => (x"c1",x"49",x"70",x"30"),
  1597 => (x"7a",x"97",x"71",x"89"),
  1598 => (x"bf",x"d0",x"f1",x"c2"),
  1599 => (x"97",x"29",x"6e",x"49"),
  1600 => (x"71",x"48",x"4a",x"6a"),
  1601 => (x"a6",x"f4",x"c0",x"98"),
  1602 => (x"48",x"66",x"c4",x"58"),
  1603 => (x"a6",x"cc",x"80",x"c4"),
  1604 => (x"bf",x"66",x"c8",x"58"),
  1605 => (x"66",x"e4",x"c0",x"4c"),
  1606 => (x"a8",x"66",x"cc",x"48"),
  1607 => (x"87",x"c5",x"c0",x"02"),
  1608 => (x"c2",x"c0",x"7e",x"c0"),
  1609 => (x"6e",x"7e",x"c1",x"87"),
  1610 => (x"1e",x"e0",x"c0",x"1e"),
  1611 => (x"d5",x"ff",x"49",x"74"),
  1612 => (x"86",x"c8",x"87",x"f6"),
  1613 => (x"b7",x"c0",x"4d",x"70"),
  1614 => (x"d4",x"c1",x"06",x"ad"),
  1615 => (x"c8",x"84",x"75",x"87"),
  1616 => (x"c0",x"49",x"bf",x"66"),
  1617 => (x"89",x"74",x"81",x"e0"),
  1618 => (x"f8",x"c9",x"c1",x"4b"),
  1619 => (x"de",x"fe",x"71",x"4a"),
  1620 => (x"84",x"c2",x"87",x"ee"),
  1621 => (x"e8",x"c0",x"7e",x"74"),
  1622 => (x"80",x"c1",x"48",x"66"),
  1623 => (x"58",x"a6",x"ec",x"c0"),
  1624 => (x"49",x"66",x"f0",x"c0"),
  1625 => (x"a9",x"70",x"81",x"c1"),
  1626 => (x"87",x"c5",x"c0",x"02"),
  1627 => (x"c2",x"c0",x"4c",x"c0"),
  1628 => (x"74",x"4c",x"c1",x"87"),
  1629 => (x"bf",x"66",x"cc",x"1e"),
  1630 => (x"81",x"e0",x"c0",x"49"),
  1631 => (x"71",x"89",x"66",x"c4"),
  1632 => (x"49",x"66",x"c8",x"1e"),
  1633 => (x"87",x"e0",x"d4",x"ff"),
  1634 => (x"b7",x"c0",x"86",x"c8"),
  1635 => (x"c5",x"ff",x"01",x"a8"),
  1636 => (x"66",x"e8",x"c0",x"87"),
  1637 => (x"87",x"d3",x"c0",x"02"),
  1638 => (x"c9",x"49",x"66",x"c4"),
  1639 => (x"66",x"e8",x"c0",x"81"),
  1640 => (x"48",x"66",x"c4",x"51"),
  1641 => (x"78",x"fa",x"d5",x"c1"),
  1642 => (x"c4",x"87",x"ce",x"c0"),
  1643 => (x"81",x"c9",x"49",x"66"),
  1644 => (x"66",x"c4",x"51",x"c2"),
  1645 => (x"f8",x"d7",x"c1",x"48"),
  1646 => (x"48",x"66",x"d4",x"78"),
  1647 => (x"04",x"a8",x"66",x"d8"),
  1648 => (x"d4",x"87",x"cb",x"c0"),
  1649 => (x"80",x"c1",x"48",x"66"),
  1650 => (x"c0",x"58",x"a6",x"d8"),
  1651 => (x"66",x"d8",x"87",x"d1"),
  1652 => (x"dc",x"88",x"c1",x"48"),
  1653 => (x"c6",x"c0",x"58",x"a6"),
  1654 => (x"f7",x"d2",x"ff",x"87"),
  1655 => (x"cc",x"4d",x"70",x"87"),
  1656 => (x"78",x"c0",x"48",x"a6"),
  1657 => (x"ff",x"87",x"c6",x"c0"),
  1658 => (x"70",x"87",x"e9",x"d2"),
  1659 => (x"66",x"e0",x"c0",x"4d"),
  1660 => (x"c0",x"80",x"c1",x"48"),
  1661 => (x"75",x"58",x"a6",x"e4"),
  1662 => (x"cb",x"c0",x"02",x"9d"),
  1663 => (x"48",x"66",x"d4",x"87"),
  1664 => (x"a8",x"66",x"cc",x"c1"),
  1665 => (x"87",x"da",x"f4",x"04"),
  1666 => (x"c7",x"48",x"66",x"d4"),
  1667 => (x"e1",x"c0",x"03",x"a8"),
  1668 => (x"4c",x"66",x"d4",x"87"),
  1669 => (x"48",x"e8",x"f2",x"c2"),
  1670 => (x"49",x"74",x"78",x"c0"),
  1671 => (x"c4",x"c1",x"91",x"cc"),
  1672 => (x"a1",x"c4",x"81",x"66"),
  1673 => (x"c0",x"4a",x"6a",x"4a"),
  1674 => (x"84",x"c1",x"79",x"52"),
  1675 => (x"ff",x"04",x"ac",x"c7"),
  1676 => (x"e4",x"c0",x"87",x"e2"),
  1677 => (x"e2",x"c0",x"02",x"66"),
  1678 => (x"66",x"c4",x"c1",x"87"),
  1679 => (x"81",x"d4",x"c1",x"49"),
  1680 => (x"4a",x"66",x"c4",x"c1"),
  1681 => (x"c0",x"82",x"dc",x"c1"),
  1682 => (x"ec",x"d4",x"c1",x"52"),
  1683 => (x"66",x"c4",x"c1",x"79"),
  1684 => (x"81",x"d8",x"c1",x"49"),
  1685 => (x"79",x"fc",x"c9",x"c1"),
  1686 => (x"c1",x"87",x"d6",x"c0"),
  1687 => (x"c1",x"49",x"66",x"c4"),
  1688 => (x"c4",x"c1",x"81",x"d4"),
  1689 => (x"d8",x"c1",x"4a",x"66"),
  1690 => (x"c4",x"ca",x"c1",x"82"),
  1691 => (x"e3",x"d4",x"c1",x"7a"),
  1692 => (x"ca",x"d8",x"c1",x"79"),
  1693 => (x"66",x"c4",x"c1",x"4a"),
  1694 => (x"81",x"e0",x"c1",x"49"),
  1695 => (x"d0",x"ff",x"79",x"72"),
  1696 => (x"66",x"d0",x"87",x"c9"),
  1697 => (x"8e",x"cc",x"ff",x"48"),
  1698 => (x"4c",x"26",x"4d",x"26"),
  1699 => (x"4f",x"26",x"4b",x"26"),
  1700 => (x"c2",x"1e",x"c7",x"1e"),
  1701 => (x"1e",x"bf",x"e4",x"f2"),
  1702 => (x"1e",x"f8",x"ec",x"c1"),
  1703 => (x"97",x"d4",x"f1",x"c2"),
  1704 => (x"f7",x"ee",x"49",x"bf"),
  1705 => (x"f8",x"ec",x"c1",x"87"),
  1706 => (x"ed",x"e1",x"c0",x"49"),
  1707 => (x"26",x"8e",x"f4",x"87"),
  1708 => (x"1e",x"73",x"1e",x"4f"),
  1709 => (x"c2",x"87",x"cf",x"c7"),
  1710 => (x"c0",x"48",x"f0",x"f2"),
  1711 => (x"48",x"d4",x"ff",x"50"),
  1712 => (x"c1",x"78",x"ff",x"c3"),
  1713 => (x"fe",x"49",x"cc",x"ca"),
  1714 => (x"fe",x"87",x"dc",x"d7"),
  1715 => (x"70",x"87",x"f1",x"e2"),
  1716 => (x"87",x"cd",x"02",x"98"),
  1717 => (x"87",x"cf",x"ec",x"fe"),
  1718 => (x"c4",x"02",x"98",x"70"),
  1719 => (x"c2",x"4a",x"c1",x"87"),
  1720 => (x"72",x"4a",x"c0",x"87"),
  1721 => (x"87",x"c8",x"02",x"9a"),
  1722 => (x"49",x"d8",x"ca",x"c1"),
  1723 => (x"87",x"f7",x"d6",x"fe"),
  1724 => (x"48",x"e4",x"f2",x"c2"),
  1725 => (x"f1",x"c2",x"78",x"c0"),
  1726 => (x"50",x"c0",x"48",x"d4"),
  1727 => (x"87",x"d0",x"fe",x"49"),
  1728 => (x"87",x"f1",x"f6",x"c0"),
  1729 => (x"02",x"9b",x"4b",x"70"),
  1730 => (x"ee",x"c1",x"87",x"cf"),
  1731 => (x"49",x"c7",x"5b",x"d4"),
  1732 => (x"c1",x"87",x"f9",x"de"),
  1733 => (x"d4",x"e0",x"c0",x"49"),
  1734 => (x"87",x"f3",x"c2",x"87"),
  1735 => (x"87",x"da",x"e1",x"c0"),
  1736 => (x"87",x"f5",x"ef",x"c0"),
  1737 => (x"26",x"87",x"f5",x"ff"),
  1738 => (x"00",x"4f",x"26",x"4b"),
  1739 => (x"00",x"00",x"00",x"00"),
  1740 => (x"00",x"00",x"00",x"00"),
  1741 => (x"00",x"00",x"00",x"01"),
  1742 => (x"00",x"00",x"11",x"d6"),
  1743 => (x"00",x"00",x"2c",x"bc"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"00",x"00",x"11",x"d6"),
  1746 => (x"00",x"00",x"2c",x"da"),
  1747 => (x"00",x"00",x"00",x"00"),
  1748 => (x"00",x"00",x"11",x"d6"),
  1749 => (x"00",x"00",x"2c",x"f8"),
  1750 => (x"00",x"00",x"00",x"00"),
  1751 => (x"00",x"00",x"11",x"d6"),
  1752 => (x"00",x"00",x"2d",x"16"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"11",x"d6"),
  1755 => (x"00",x"00",x"2d",x"34"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"11",x"d6"),
  1758 => (x"00",x"00",x"2d",x"52"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"11",x"d6"),
  1761 => (x"00",x"00",x"2d",x"70"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"15",x"2c"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"12",x"d0"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"12",x"9c"),
  1770 => (x"db",x"86",x"fc",x"1e"),
  1771 => (x"fc",x"7e",x"70",x"87"),
  1772 => (x"1e",x"4f",x"26",x"8e"),
  1773 => (x"c0",x"48",x"f0",x"fe"),
  1774 => (x"79",x"09",x"cd",x"78"),
  1775 => (x"1e",x"4f",x"26",x"09"),
  1776 => (x"49",x"e8",x"ee",x"c1"),
  1777 => (x"4f",x"26",x"87",x"ed"),
  1778 => (x"bf",x"f0",x"fe",x"1e"),
  1779 => (x"1e",x"4f",x"26",x"48"),
  1780 => (x"c1",x"48",x"f0",x"fe"),
  1781 => (x"1e",x"4f",x"26",x"78"),
  1782 => (x"c0",x"48",x"f0",x"fe"),
  1783 => (x"1e",x"4f",x"26",x"78"),
  1784 => (x"52",x"c0",x"4a",x"71"),
  1785 => (x"0e",x"4f",x"26",x"51"),
  1786 => (x"5d",x"5c",x"5b",x"5e"),
  1787 => (x"71",x"86",x"f4",x"0e"),
  1788 => (x"7e",x"6d",x"97",x"4d"),
  1789 => (x"97",x"4c",x"a5",x"c1"),
  1790 => (x"a6",x"c8",x"48",x"6c"),
  1791 => (x"c4",x"48",x"6e",x"58"),
  1792 => (x"c5",x"05",x"a8",x"66"),
  1793 => (x"c0",x"48",x"ff",x"87"),
  1794 => (x"ca",x"ff",x"87",x"e6"),
  1795 => (x"49",x"a5",x"c2",x"87"),
  1796 => (x"71",x"4b",x"6c",x"97"),
  1797 => (x"6b",x"97",x"4b",x"a3"),
  1798 => (x"7e",x"6c",x"97",x"4b"),
  1799 => (x"80",x"c1",x"48",x"6e"),
  1800 => (x"c7",x"58",x"a6",x"c8"),
  1801 => (x"58",x"a6",x"cc",x"98"),
  1802 => (x"fe",x"7c",x"97",x"70"),
  1803 => (x"48",x"73",x"87",x"e1"),
  1804 => (x"4d",x"26",x"8e",x"f4"),
  1805 => (x"4b",x"26",x"4c",x"26"),
  1806 => (x"73",x"1e",x"4f",x"26"),
  1807 => (x"fe",x"86",x"f4",x"1e"),
  1808 => (x"bf",x"e0",x"87",x"d5"),
  1809 => (x"e0",x"c0",x"49",x"4b"),
  1810 => (x"c0",x"02",x"99",x"c0"),
  1811 => (x"4a",x"73",x"87",x"ea"),
  1812 => (x"c2",x"9a",x"ff",x"c3"),
  1813 => (x"bf",x"97",x"e4",x"f6"),
  1814 => (x"e6",x"f6",x"c2",x"49"),
  1815 => (x"c2",x"51",x"72",x"81"),
  1816 => (x"bf",x"97",x"e4",x"f6"),
  1817 => (x"c1",x"48",x"6e",x"7e"),
  1818 => (x"58",x"a6",x"c8",x"80"),
  1819 => (x"a6",x"cc",x"98",x"c7"),
  1820 => (x"e4",x"f6",x"c2",x"58"),
  1821 => (x"50",x"66",x"c8",x"48"),
  1822 => (x"70",x"87",x"cd",x"fd"),
  1823 => (x"87",x"cf",x"fd",x"7e"),
  1824 => (x"4b",x"26",x"8e",x"f4"),
  1825 => (x"c2",x"1e",x"4f",x"26"),
  1826 => (x"fd",x"49",x"e4",x"f6"),
  1827 => (x"f0",x"c1",x"87",x"d1"),
  1828 => (x"de",x"fc",x"49",x"fa"),
  1829 => (x"87",x"e8",x"c4",x"87"),
  1830 => (x"5e",x"0e",x"4f",x"26"),
  1831 => (x"0e",x"5d",x"5c",x"5b"),
  1832 => (x"7e",x"71",x"86",x"fc"),
  1833 => (x"c2",x"4d",x"d4",x"ff"),
  1834 => (x"fc",x"49",x"e4",x"f6"),
  1835 => (x"4b",x"70",x"87",x"f9"),
  1836 => (x"04",x"ab",x"b7",x"c0"),
  1837 => (x"c3",x"87",x"f5",x"c2"),
  1838 => (x"c9",x"05",x"ab",x"f0"),
  1839 => (x"f8",x"f5",x"c1",x"87"),
  1840 => (x"c2",x"78",x"c1",x"48"),
  1841 => (x"e0",x"c3",x"87",x"d6"),
  1842 => (x"87",x"c9",x"05",x"ab"),
  1843 => (x"48",x"fc",x"f5",x"c1"),
  1844 => (x"c7",x"c2",x"78",x"c1"),
  1845 => (x"fc",x"f5",x"c1",x"87"),
  1846 => (x"87",x"c6",x"02",x"bf"),
  1847 => (x"4c",x"a3",x"c0",x"c2"),
  1848 => (x"4c",x"73",x"87",x"c2"),
  1849 => (x"bf",x"f8",x"f5",x"c1"),
  1850 => (x"87",x"e0",x"c0",x"02"),
  1851 => (x"b7",x"c4",x"49",x"74"),
  1852 => (x"f6",x"c1",x"91",x"29"),
  1853 => (x"4a",x"74",x"81",x"c0"),
  1854 => (x"92",x"c2",x"9a",x"cf"),
  1855 => (x"30",x"72",x"48",x"c1"),
  1856 => (x"ba",x"ff",x"4a",x"70"),
  1857 => (x"98",x"69",x"48",x"72"),
  1858 => (x"87",x"db",x"79",x"70"),
  1859 => (x"b7",x"c4",x"49",x"74"),
  1860 => (x"f6",x"c1",x"91",x"29"),
  1861 => (x"4a",x"74",x"81",x"c0"),
  1862 => (x"92",x"c2",x"9a",x"cf"),
  1863 => (x"30",x"72",x"48",x"c3"),
  1864 => (x"69",x"48",x"4a",x"70"),
  1865 => (x"6e",x"79",x"70",x"b0"),
  1866 => (x"87",x"e4",x"c0",x"05"),
  1867 => (x"c8",x"48",x"d0",x"ff"),
  1868 => (x"7d",x"c5",x"78",x"e1"),
  1869 => (x"bf",x"fc",x"f5",x"c1"),
  1870 => (x"c3",x"87",x"c3",x"02"),
  1871 => (x"f5",x"c1",x"7d",x"e0"),
  1872 => (x"c3",x"02",x"bf",x"f8"),
  1873 => (x"7d",x"f0",x"c3",x"87"),
  1874 => (x"d0",x"ff",x"7d",x"73"),
  1875 => (x"78",x"e0",x"c0",x"48"),
  1876 => (x"48",x"fc",x"f5",x"c1"),
  1877 => (x"f5",x"c1",x"78",x"c0"),
  1878 => (x"78",x"c0",x"48",x"f8"),
  1879 => (x"49",x"e4",x"f6",x"c2"),
  1880 => (x"70",x"87",x"c4",x"fa"),
  1881 => (x"ab",x"b7",x"c0",x"4b"),
  1882 => (x"87",x"cb",x"fd",x"03"),
  1883 => (x"8e",x"fc",x"48",x"c0"),
  1884 => (x"4c",x"26",x"4d",x"26"),
  1885 => (x"4f",x"26",x"4b",x"26"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"00",x"00",x"00",x"00"),
  1894 => (x"00",x"00",x"00",x"00"),
  1895 => (x"00",x"00",x"00",x"00"),
  1896 => (x"00",x"00",x"00",x"00"),
  1897 => (x"00",x"00",x"00",x"00"),
  1898 => (x"00",x"00",x"00",x"00"),
  1899 => (x"00",x"00",x"00",x"00"),
  1900 => (x"00",x"00",x"00",x"00"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"00",x"00",x"00",x"00"),
  1904 => (x"72",x"4a",x"c0",x"1e"),
  1905 => (x"c1",x"91",x"c4",x"49"),
  1906 => (x"c0",x"81",x"c0",x"f6"),
  1907 => (x"d0",x"82",x"c1",x"79"),
  1908 => (x"ee",x"04",x"aa",x"b7"),
  1909 => (x"0e",x"4f",x"26",x"87"),
  1910 => (x"5d",x"5c",x"5b",x"5e"),
  1911 => (x"f7",x"4d",x"71",x"0e"),
  1912 => (x"4a",x"75",x"87",x"f5"),
  1913 => (x"92",x"2a",x"b7",x"c4"),
  1914 => (x"82",x"c0",x"f6",x"c1"),
  1915 => (x"9c",x"cf",x"4c",x"75"),
  1916 => (x"49",x"6a",x"94",x"c2"),
  1917 => (x"c3",x"2b",x"74",x"4b"),
  1918 => (x"74",x"48",x"c2",x"9b"),
  1919 => (x"ff",x"4c",x"70",x"30"),
  1920 => (x"71",x"48",x"74",x"bc"),
  1921 => (x"f7",x"7a",x"70",x"98"),
  1922 => (x"48",x"73",x"87",x"c5"),
  1923 => (x"4c",x"26",x"4d",x"26"),
  1924 => (x"4f",x"26",x"4b",x"26"),
  1925 => (x"48",x"d0",x"ff",x"1e"),
  1926 => (x"71",x"78",x"e1",x"c8"),
  1927 => (x"08",x"d4",x"ff",x"48"),
  1928 => (x"1e",x"4f",x"26",x"78"),
  1929 => (x"c8",x"48",x"d0",x"ff"),
  1930 => (x"48",x"71",x"78",x"e1"),
  1931 => (x"78",x"08",x"d4",x"ff"),
  1932 => (x"ff",x"48",x"66",x"c4"),
  1933 => (x"26",x"78",x"08",x"d4"),
  1934 => (x"4a",x"71",x"1e",x"4f"),
  1935 => (x"1e",x"49",x"66",x"c4"),
  1936 => (x"de",x"ff",x"49",x"72"),
  1937 => (x"48",x"d0",x"ff",x"87"),
  1938 => (x"fc",x"78",x"e0",x"c0"),
  1939 => (x"1e",x"4f",x"26",x"8e"),
  1940 => (x"4a",x"71",x"1e",x"73"),
  1941 => (x"ab",x"b7",x"c2",x"4b"),
  1942 => (x"a3",x"87",x"c8",x"03"),
  1943 => (x"ff",x"c3",x"4a",x"49"),
  1944 => (x"ce",x"87",x"c7",x"9a"),
  1945 => (x"c3",x"4a",x"49",x"a3"),
  1946 => (x"66",x"c8",x"9a",x"ff"),
  1947 => (x"49",x"72",x"1e",x"49"),
  1948 => (x"fc",x"87",x"c6",x"ff"),
  1949 => (x"26",x"4b",x"26",x"8e"),
  1950 => (x"d0",x"ff",x"1e",x"4f"),
  1951 => (x"78",x"c9",x"c8",x"48"),
  1952 => (x"d4",x"ff",x"48",x"71"),
  1953 => (x"4f",x"26",x"78",x"08"),
  1954 => (x"49",x"4a",x"71",x"1e"),
  1955 => (x"d0",x"ff",x"87",x"eb"),
  1956 => (x"26",x"78",x"c8",x"48"),
  1957 => (x"1e",x"73",x"1e",x"4f"),
  1958 => (x"f6",x"c2",x"4b",x"71"),
  1959 => (x"c3",x"02",x"bf",x"fc"),
  1960 => (x"87",x"eb",x"c2",x"87"),
  1961 => (x"c8",x"48",x"d0",x"ff"),
  1962 => (x"48",x"73",x"78",x"c9"),
  1963 => (x"ff",x"b0",x"e0",x"c0"),
  1964 => (x"c2",x"78",x"08",x"d4"),
  1965 => (x"c0",x"48",x"f0",x"f6"),
  1966 => (x"02",x"66",x"c8",x"78"),
  1967 => (x"ff",x"c3",x"87",x"c5"),
  1968 => (x"c0",x"87",x"c2",x"49"),
  1969 => (x"f8",x"f6",x"c2",x"49"),
  1970 => (x"02",x"66",x"cc",x"59"),
  1971 => (x"d5",x"c5",x"87",x"c6"),
  1972 => (x"87",x"c4",x"4a",x"d5"),
  1973 => (x"4a",x"ff",x"ff",x"cf"),
  1974 => (x"5a",x"fc",x"f6",x"c2"),
  1975 => (x"48",x"fc",x"f6",x"c2"),
  1976 => (x"4b",x"26",x"78",x"c1"),
  1977 => (x"5e",x"0e",x"4f",x"26"),
  1978 => (x"0e",x"5d",x"5c",x"5b"),
  1979 => (x"f6",x"c2",x"4d",x"71"),
  1980 => (x"75",x"4b",x"bf",x"f8"),
  1981 => (x"87",x"cb",x"02",x"9d"),
  1982 => (x"c1",x"91",x"c8",x"49"),
  1983 => (x"71",x"4a",x"cc",x"fa"),
  1984 => (x"c1",x"87",x"c4",x"82"),
  1985 => (x"c0",x"4a",x"cc",x"fe"),
  1986 => (x"73",x"49",x"12",x"4c"),
  1987 => (x"f4",x"f6",x"c2",x"99"),
  1988 => (x"b8",x"71",x"48",x"bf"),
  1989 => (x"78",x"08",x"d4",x"ff"),
  1990 => (x"84",x"2b",x"b7",x"c1"),
  1991 => (x"04",x"ac",x"b7",x"c8"),
  1992 => (x"f6",x"c2",x"87",x"e7"),
  1993 => (x"c8",x"48",x"bf",x"f0"),
  1994 => (x"f4",x"f6",x"c2",x"80"),
  1995 => (x"26",x"4d",x"26",x"58"),
  1996 => (x"26",x"4b",x"26",x"4c"),
  1997 => (x"1e",x"73",x"1e",x"4f"),
  1998 => (x"4a",x"13",x"4b",x"71"),
  1999 => (x"87",x"cb",x"02",x"9a"),
  2000 => (x"e1",x"fe",x"49",x"72"),
  2001 => (x"9a",x"4a",x"13",x"87"),
  2002 => (x"26",x"87",x"f5",x"05"),
  2003 => (x"1e",x"4f",x"26",x"4b"),
  2004 => (x"bf",x"f0",x"f6",x"c2"),
  2005 => (x"f0",x"f6",x"c2",x"49"),
  2006 => (x"78",x"a1",x"c1",x"48"),
  2007 => (x"a9",x"b7",x"c0",x"c4"),
  2008 => (x"ff",x"87",x"db",x"03"),
  2009 => (x"f6",x"c2",x"48",x"d4"),
  2010 => (x"c2",x"78",x"bf",x"f4"),
  2011 => (x"49",x"bf",x"f0",x"f6"),
  2012 => (x"48",x"f0",x"f6",x"c2"),
  2013 => (x"c4",x"78",x"a1",x"c1"),
  2014 => (x"04",x"a9",x"b7",x"c0"),
  2015 => (x"d0",x"ff",x"87",x"e5"),
  2016 => (x"c2",x"78",x"c8",x"48"),
  2017 => (x"c0",x"48",x"fc",x"f6"),
  2018 => (x"00",x"4f",x"26",x"78"),
  2019 => (x"00",x"00",x"00",x"00"),
  2020 => (x"00",x"00",x"00",x"00"),
  2021 => (x"5f",x"00",x"00",x"00"),
  2022 => (x"00",x"00",x"00",x"5f"),
  2023 => (x"00",x"03",x"03",x"00"),
  2024 => (x"00",x"00",x"03",x"03"),
  2025 => (x"14",x"7f",x"7f",x"14"),
  2026 => (x"00",x"14",x"7f",x"7f"),
  2027 => (x"6b",x"2e",x"24",x"00"),
  2028 => (x"00",x"12",x"3a",x"6b"),
  2029 => (x"18",x"36",x"6a",x"4c"),
  2030 => (x"00",x"32",x"56",x"6c"),
  2031 => (x"59",x"4f",x"7e",x"30"),
  2032 => (x"40",x"68",x"3a",x"77"),
  2033 => (x"07",x"04",x"00",x"00"),
  2034 => (x"00",x"00",x"00",x"03"),
  2035 => (x"3e",x"1c",x"00",x"00"),
  2036 => (x"00",x"00",x"41",x"63"),
  2037 => (x"63",x"41",x"00",x"00"),
  2038 => (x"00",x"00",x"1c",x"3e"),
  2039 => (x"1c",x"3e",x"2a",x"08"),
  2040 => (x"08",x"2a",x"3e",x"1c"),
  2041 => (x"3e",x"08",x"08",x"00"),
  2042 => (x"00",x"08",x"08",x"3e"),
  2043 => (x"e0",x"80",x"00",x"00"),
  2044 => (x"00",x"00",x"00",x"60"),
  2045 => (x"08",x"08",x"08",x"00"),
  2046 => (x"00",x"08",x"08",x"08"),
  2047 => (x"60",x"00",x"00",x"00"),
  2048 => (x"00",x"00",x"00",x"60"),
  2049 => (x"18",x"30",x"60",x"40"),
  2050 => (x"01",x"03",x"06",x"0c"),
  2051 => (x"59",x"7f",x"3e",x"00"),
  2052 => (x"00",x"3e",x"7f",x"4d"),
  2053 => (x"7f",x"06",x"04",x"00"),
  2054 => (x"00",x"00",x"00",x"7f"),
  2055 => (x"71",x"63",x"42",x"00"),
  2056 => (x"00",x"46",x"4f",x"59"),
  2057 => (x"49",x"63",x"22",x"00"),
  2058 => (x"00",x"36",x"7f",x"49"),
  2059 => (x"13",x"16",x"1c",x"18"),
  2060 => (x"00",x"10",x"7f",x"7f"),
  2061 => (x"45",x"67",x"27",x"00"),
  2062 => (x"00",x"39",x"7d",x"45"),
  2063 => (x"4b",x"7e",x"3c",x"00"),
  2064 => (x"00",x"30",x"79",x"49"),
  2065 => (x"71",x"01",x"01",x"00"),
  2066 => (x"00",x"07",x"0f",x"79"),
  2067 => (x"49",x"7f",x"36",x"00"),
  2068 => (x"00",x"36",x"7f",x"49"),
  2069 => (x"49",x"4f",x"06",x"00"),
  2070 => (x"00",x"1e",x"3f",x"69"),
  2071 => (x"66",x"00",x"00",x"00"),
  2072 => (x"00",x"00",x"00",x"66"),
  2073 => (x"e6",x"80",x"00",x"00"),
  2074 => (x"00",x"00",x"00",x"66"),
  2075 => (x"14",x"08",x"08",x"00"),
  2076 => (x"00",x"22",x"22",x"14"),
  2077 => (x"14",x"14",x"14",x"00"),
  2078 => (x"00",x"14",x"14",x"14"),
  2079 => (x"14",x"22",x"22",x"00"),
  2080 => (x"00",x"08",x"08",x"14"),
  2081 => (x"51",x"03",x"02",x"00"),
  2082 => (x"00",x"06",x"0f",x"59"),
  2083 => (x"5d",x"41",x"7f",x"3e"),
  2084 => (x"00",x"1e",x"1f",x"55"),
  2085 => (x"09",x"7f",x"7e",x"00"),
  2086 => (x"00",x"7e",x"7f",x"09"),
  2087 => (x"49",x"7f",x"7f",x"00"),
  2088 => (x"00",x"36",x"7f",x"49"),
  2089 => (x"63",x"3e",x"1c",x"00"),
  2090 => (x"00",x"41",x"41",x"41"),
  2091 => (x"41",x"7f",x"7f",x"00"),
  2092 => (x"00",x"1c",x"3e",x"63"),
  2093 => (x"49",x"7f",x"7f",x"00"),
  2094 => (x"00",x"41",x"41",x"49"),
  2095 => (x"09",x"7f",x"7f",x"00"),
  2096 => (x"00",x"01",x"01",x"09"),
  2097 => (x"41",x"7f",x"3e",x"00"),
  2098 => (x"00",x"7a",x"7b",x"49"),
  2099 => (x"08",x"7f",x"7f",x"00"),
  2100 => (x"00",x"7f",x"7f",x"08"),
  2101 => (x"7f",x"41",x"00",x"00"),
  2102 => (x"00",x"00",x"41",x"7f"),
  2103 => (x"40",x"60",x"20",x"00"),
  2104 => (x"00",x"3f",x"7f",x"40"),
  2105 => (x"1c",x"08",x"7f",x"7f"),
  2106 => (x"00",x"41",x"63",x"36"),
  2107 => (x"40",x"7f",x"7f",x"00"),
  2108 => (x"00",x"40",x"40",x"40"),
  2109 => (x"0c",x"06",x"7f",x"7f"),
  2110 => (x"00",x"7f",x"7f",x"06"),
  2111 => (x"0c",x"06",x"7f",x"7f"),
  2112 => (x"00",x"7f",x"7f",x"18"),
  2113 => (x"41",x"7f",x"3e",x"00"),
  2114 => (x"00",x"3e",x"7f",x"41"),
  2115 => (x"09",x"7f",x"7f",x"00"),
  2116 => (x"00",x"06",x"0f",x"09"),
  2117 => (x"61",x"41",x"7f",x"3e"),
  2118 => (x"00",x"40",x"7e",x"7f"),
  2119 => (x"09",x"7f",x"7f",x"00"),
  2120 => (x"00",x"66",x"7f",x"19"),
  2121 => (x"4d",x"6f",x"26",x"00"),
  2122 => (x"00",x"32",x"7b",x"59"),
  2123 => (x"7f",x"01",x"01",x"00"),
  2124 => (x"00",x"01",x"01",x"7f"),
  2125 => (x"40",x"7f",x"3f",x"00"),
  2126 => (x"00",x"3f",x"7f",x"40"),
  2127 => (x"70",x"3f",x"0f",x"00"),
  2128 => (x"00",x"0f",x"3f",x"70"),
  2129 => (x"18",x"30",x"7f",x"7f"),
  2130 => (x"00",x"7f",x"7f",x"30"),
  2131 => (x"1c",x"36",x"63",x"41"),
  2132 => (x"41",x"63",x"36",x"1c"),
  2133 => (x"7c",x"06",x"03",x"01"),
  2134 => (x"01",x"03",x"06",x"7c"),
  2135 => (x"4d",x"59",x"71",x"61"),
  2136 => (x"00",x"41",x"43",x"47"),
  2137 => (x"7f",x"7f",x"00",x"00"),
  2138 => (x"00",x"00",x"41",x"41"),
  2139 => (x"0c",x"06",x"03",x"01"),
  2140 => (x"40",x"60",x"30",x"18"),
  2141 => (x"41",x"41",x"00",x"00"),
  2142 => (x"00",x"00",x"7f",x"7f"),
  2143 => (x"03",x"06",x"0c",x"08"),
  2144 => (x"00",x"08",x"0c",x"06"),
  2145 => (x"80",x"80",x"80",x"80"),
  2146 => (x"00",x"80",x"80",x"80"),
  2147 => (x"03",x"00",x"00",x"00"),
  2148 => (x"00",x"00",x"04",x"07"),
  2149 => (x"54",x"74",x"20",x"00"),
  2150 => (x"00",x"78",x"7c",x"54"),
  2151 => (x"44",x"7f",x"7f",x"00"),
  2152 => (x"00",x"38",x"7c",x"44"),
  2153 => (x"44",x"7c",x"38",x"00"),
  2154 => (x"00",x"00",x"44",x"44"),
  2155 => (x"44",x"7c",x"38",x"00"),
  2156 => (x"00",x"7f",x"7f",x"44"),
  2157 => (x"54",x"7c",x"38",x"00"),
  2158 => (x"00",x"18",x"5c",x"54"),
  2159 => (x"7f",x"7e",x"04",x"00"),
  2160 => (x"00",x"00",x"05",x"05"),
  2161 => (x"a4",x"bc",x"18",x"00"),
  2162 => (x"00",x"7c",x"fc",x"a4"),
  2163 => (x"04",x"7f",x"7f",x"00"),
  2164 => (x"00",x"78",x"7c",x"04"),
  2165 => (x"3d",x"00",x"00",x"00"),
  2166 => (x"00",x"00",x"40",x"7d"),
  2167 => (x"80",x"80",x"80",x"00"),
  2168 => (x"00",x"00",x"7d",x"fd"),
  2169 => (x"10",x"7f",x"7f",x"00"),
  2170 => (x"00",x"44",x"6c",x"38"),
  2171 => (x"3f",x"00",x"00",x"00"),
  2172 => (x"00",x"00",x"40",x"7f"),
  2173 => (x"18",x"0c",x"7c",x"7c"),
  2174 => (x"00",x"78",x"7c",x"0c"),
  2175 => (x"04",x"7c",x"7c",x"00"),
  2176 => (x"00",x"78",x"7c",x"04"),
  2177 => (x"44",x"7c",x"38",x"00"),
  2178 => (x"00",x"38",x"7c",x"44"),
  2179 => (x"24",x"fc",x"fc",x"00"),
  2180 => (x"00",x"18",x"3c",x"24"),
  2181 => (x"24",x"3c",x"18",x"00"),
  2182 => (x"00",x"fc",x"fc",x"24"),
  2183 => (x"04",x"7c",x"7c",x"00"),
  2184 => (x"00",x"08",x"0c",x"04"),
  2185 => (x"54",x"5c",x"48",x"00"),
  2186 => (x"00",x"20",x"74",x"54"),
  2187 => (x"7f",x"3f",x"04",x"00"),
  2188 => (x"00",x"00",x"44",x"44"),
  2189 => (x"40",x"7c",x"3c",x"00"),
  2190 => (x"00",x"7c",x"7c",x"40"),
  2191 => (x"60",x"3c",x"1c",x"00"),
  2192 => (x"00",x"1c",x"3c",x"60"),
  2193 => (x"30",x"60",x"7c",x"3c"),
  2194 => (x"00",x"3c",x"7c",x"60"),
  2195 => (x"10",x"38",x"6c",x"44"),
  2196 => (x"00",x"44",x"6c",x"38"),
  2197 => (x"e0",x"bc",x"1c",x"00"),
  2198 => (x"00",x"1c",x"3c",x"60"),
  2199 => (x"74",x"64",x"44",x"00"),
  2200 => (x"00",x"44",x"4c",x"5c"),
  2201 => (x"3e",x"08",x"08",x"00"),
  2202 => (x"00",x"41",x"41",x"77"),
  2203 => (x"7f",x"00",x"00",x"00"),
  2204 => (x"00",x"00",x"00",x"7f"),
  2205 => (x"77",x"41",x"41",x"00"),
  2206 => (x"00",x"08",x"08",x"3e"),
  2207 => (x"03",x"01",x"01",x"02"),
  2208 => (x"00",x"01",x"02",x"02"),
  2209 => (x"7f",x"7f",x"7f",x"7f"),
  2210 => (x"00",x"7f",x"7f",x"7f"),
  2211 => (x"1c",x"1c",x"08",x"08"),
  2212 => (x"7f",x"7f",x"3e",x"3e"),
  2213 => (x"3e",x"3e",x"7f",x"7f"),
  2214 => (x"08",x"08",x"1c",x"1c"),
  2215 => (x"7c",x"18",x"10",x"00"),
  2216 => (x"00",x"10",x"18",x"7c"),
  2217 => (x"7c",x"30",x"10",x"00"),
  2218 => (x"00",x"10",x"30",x"7c"),
  2219 => (x"60",x"60",x"30",x"10"),
  2220 => (x"00",x"06",x"1e",x"78"),
  2221 => (x"18",x"3c",x"66",x"42"),
  2222 => (x"00",x"42",x"66",x"3c"),
  2223 => (x"c2",x"6a",x"38",x"78"),
  2224 => (x"00",x"38",x"6c",x"c6"),
  2225 => (x"60",x"00",x"00",x"60"),
  2226 => (x"00",x"60",x"00",x"00"),
  2227 => (x"5c",x"5b",x"5e",x"0e"),
  2228 => (x"86",x"fc",x"0e",x"5d"),
  2229 => (x"f7",x"c2",x"7e",x"71"),
  2230 => (x"c0",x"4c",x"bf",x"c4"),
  2231 => (x"c4",x"1e",x"c0",x"4b"),
  2232 => (x"c4",x"02",x"ab",x"66"),
  2233 => (x"c2",x"4d",x"c0",x"87"),
  2234 => (x"75",x"4d",x"c1",x"87"),
  2235 => (x"ee",x"49",x"73",x"1e"),
  2236 => (x"86",x"c8",x"87",x"e3"),
  2237 => (x"ef",x"49",x"e0",x"c0"),
  2238 => (x"a4",x"c4",x"87",x"ec"),
  2239 => (x"f0",x"49",x"6a",x"4a"),
  2240 => (x"ca",x"f1",x"87",x"f3"),
  2241 => (x"c1",x"84",x"cc",x"87"),
  2242 => (x"ab",x"b7",x"c8",x"83"),
  2243 => (x"87",x"cd",x"ff",x"04"),
  2244 => (x"4d",x"26",x"8e",x"fc"),
  2245 => (x"4b",x"26",x"4c",x"26"),
  2246 => (x"71",x"1e",x"4f",x"26"),
  2247 => (x"c8",x"f7",x"c2",x"4a"),
  2248 => (x"c8",x"f7",x"c2",x"5a"),
  2249 => (x"49",x"78",x"c7",x"48"),
  2250 => (x"26",x"87",x"e1",x"fe"),
  2251 => (x"1e",x"73",x"1e",x"4f"),
  2252 => (x"0b",x"fc",x"4b",x"71"),
  2253 => (x"4a",x"73",x"0b",x"7b"),
  2254 => (x"c0",x"c1",x"9a",x"c1"),
  2255 => (x"c7",x"ed",x"49",x"a2"),
  2256 => (x"c0",x"da",x"c2",x"87"),
  2257 => (x"26",x"4b",x"26",x"5b"),
  2258 => (x"4a",x"71",x"1e",x"4f"),
  2259 => (x"72",x"1e",x"66",x"c4"),
  2260 => (x"87",x"fb",x"eb",x"49"),
  2261 => (x"4f",x"26",x"8e",x"fc"),
  2262 => (x"48",x"d4",x"ff",x"1e"),
  2263 => (x"ff",x"78",x"ff",x"c3"),
  2264 => (x"e1",x"c0",x"48",x"d0"),
  2265 => (x"48",x"d4",x"ff",x"78"),
  2266 => (x"48",x"71",x"78",x"c1"),
  2267 => (x"d4",x"ff",x"30",x"c4"),
  2268 => (x"d0",x"ff",x"78",x"08"),
  2269 => (x"78",x"e0",x"c0",x"48"),
  2270 => (x"5e",x"0e",x"4f",x"26"),
  2271 => (x"0e",x"5d",x"5c",x"5b"),
  2272 => (x"7e",x"c0",x"86",x"f4"),
  2273 => (x"ec",x"48",x"a6",x"c8"),
  2274 => (x"80",x"fc",x"78",x"bf"),
  2275 => (x"bf",x"c4",x"f7",x"c2"),
  2276 => (x"cc",x"f7",x"c2",x"78"),
  2277 => (x"bf",x"e8",x"4c",x"bf"),
  2278 => (x"fc",x"d9",x"c2",x"4d"),
  2279 => (x"f9",x"e3",x"49",x"bf"),
  2280 => (x"e8",x"49",x"c7",x"87"),
  2281 => (x"49",x"70",x"87",x"f1"),
  2282 => (x"d0",x"05",x"99",x"c2"),
  2283 => (x"f4",x"d9",x"c2",x"87"),
  2284 => (x"b9",x"ff",x"49",x"bf"),
  2285 => (x"c1",x"99",x"66",x"c8"),
  2286 => (x"f9",x"c1",x"02",x"99"),
  2287 => (x"49",x"e8",x"cf",x"87"),
  2288 => (x"70",x"87",x"fd",x"ca"),
  2289 => (x"e8",x"49",x"c7",x"4b"),
  2290 => (x"98",x"70",x"87",x"cd"),
  2291 => (x"c8",x"87",x"c9",x"05"),
  2292 => (x"99",x"c1",x"49",x"66"),
  2293 => (x"87",x"fe",x"c0",x"02"),
  2294 => (x"ec",x"48",x"a6",x"c8"),
  2295 => (x"f9",x"e2",x"78",x"bf"),
  2296 => (x"ca",x"49",x"73",x"87"),
  2297 => (x"98",x"70",x"87",x"e6"),
  2298 => (x"c2",x"87",x"d7",x"02"),
  2299 => (x"49",x"bf",x"f0",x"d9"),
  2300 => (x"d9",x"c2",x"b9",x"c1"),
  2301 => (x"fd",x"71",x"59",x"f4"),
  2302 => (x"e8",x"cf",x"87",x"de"),
  2303 => (x"87",x"c0",x"ca",x"49"),
  2304 => (x"49",x"c7",x"4b",x"70"),
  2305 => (x"70",x"87",x"d0",x"e7"),
  2306 => (x"cb",x"ff",x"05",x"98"),
  2307 => (x"49",x"66",x"c8",x"87"),
  2308 => (x"ff",x"05",x"99",x"c1"),
  2309 => (x"d9",x"c2",x"87",x"c2"),
  2310 => (x"c1",x"4a",x"bf",x"fc"),
  2311 => (x"c0",x"da",x"c2",x"ba"),
  2312 => (x"7a",x"0a",x"fc",x"5a"),
  2313 => (x"c1",x"9a",x"c1",x"0a"),
  2314 => (x"e9",x"49",x"a2",x"c0"),
  2315 => (x"da",x"c1",x"87",x"da"),
  2316 => (x"87",x"e3",x"e6",x"49"),
  2317 => (x"d9",x"c2",x"7e",x"c1"),
  2318 => (x"66",x"c8",x"48",x"f4"),
  2319 => (x"fc",x"d9",x"c2",x"78"),
  2320 => (x"e9",x"c0",x"05",x"bf"),
  2321 => (x"c3",x"49",x"75",x"87"),
  2322 => (x"1e",x"71",x"99",x"ff"),
  2323 => (x"f8",x"fb",x"49",x"c0"),
  2324 => (x"c8",x"49",x"75",x"87"),
  2325 => (x"1e",x"71",x"29",x"b7"),
  2326 => (x"ec",x"fb",x"49",x"c1"),
  2327 => (x"c3",x"86",x"c8",x"87"),
  2328 => (x"f2",x"e5",x"49",x"fd"),
  2329 => (x"49",x"fa",x"c3",x"87"),
  2330 => (x"c7",x"87",x"ec",x"e5"),
  2331 => (x"49",x"75",x"87",x"f4"),
  2332 => (x"c8",x"99",x"ff",x"c3"),
  2333 => (x"b5",x"71",x"2d",x"b7"),
  2334 => (x"c0",x"02",x"9d",x"75"),
  2335 => (x"a6",x"c8",x"87",x"e4"),
  2336 => (x"bf",x"c8",x"ff",x"48"),
  2337 => (x"49",x"66",x"c8",x"78"),
  2338 => (x"bf",x"f8",x"d9",x"c2"),
  2339 => (x"a9",x"e0",x"c2",x"89"),
  2340 => (x"87",x"c4",x"c0",x"03"),
  2341 => (x"87",x"d0",x"4d",x"c0"),
  2342 => (x"48",x"f8",x"d9",x"c2"),
  2343 => (x"c0",x"78",x"66",x"c8"),
  2344 => (x"d9",x"c2",x"87",x"c6"),
  2345 => (x"78",x"c0",x"48",x"f8"),
  2346 => (x"99",x"c8",x"49",x"75"),
  2347 => (x"87",x"ce",x"c0",x"05"),
  2348 => (x"e4",x"49",x"f5",x"c3"),
  2349 => (x"49",x"70",x"87",x"e1"),
  2350 => (x"c0",x"02",x"99",x"c2"),
  2351 => (x"f7",x"c2",x"87",x"e7"),
  2352 => (x"c0",x"02",x"bf",x"c8"),
  2353 => (x"c1",x"48",x"87",x"ca"),
  2354 => (x"cc",x"f7",x"c2",x"88"),
  2355 => (x"87",x"d3",x"c0",x"58"),
  2356 => (x"c1",x"48",x"66",x"c4"),
  2357 => (x"7e",x"70",x"80",x"e0"),
  2358 => (x"c0",x"02",x"bf",x"6e"),
  2359 => (x"ff",x"4b",x"87",x"c5"),
  2360 => (x"c1",x"0f",x"73",x"49"),
  2361 => (x"c4",x"49",x"75",x"7e"),
  2362 => (x"ce",x"c0",x"05",x"99"),
  2363 => (x"49",x"f2",x"c3",x"87"),
  2364 => (x"70",x"87",x"e4",x"e3"),
  2365 => (x"02",x"99",x"c2",x"49"),
  2366 => (x"c2",x"87",x"ea",x"c0"),
  2367 => (x"7e",x"bf",x"c8",x"f7"),
  2368 => (x"a8",x"b7",x"c7",x"48"),
  2369 => (x"87",x"cb",x"c0",x"03"),
  2370 => (x"80",x"c1",x"48",x"6e"),
  2371 => (x"58",x"cc",x"f7",x"c2"),
  2372 => (x"c4",x"87",x"d0",x"c0"),
  2373 => (x"e0",x"c1",x"4a",x"66"),
  2374 => (x"c0",x"02",x"6a",x"82"),
  2375 => (x"fe",x"4b",x"87",x"c5"),
  2376 => (x"c1",x"0f",x"73",x"49"),
  2377 => (x"49",x"fd",x"c3",x"7e"),
  2378 => (x"70",x"87",x"ec",x"e2"),
  2379 => (x"02",x"99",x"c2",x"49"),
  2380 => (x"c2",x"87",x"e6",x"c0"),
  2381 => (x"02",x"bf",x"c8",x"f7"),
  2382 => (x"c2",x"87",x"c9",x"c0"),
  2383 => (x"c0",x"48",x"c8",x"f7"),
  2384 => (x"87",x"d3",x"c0",x"78"),
  2385 => (x"c1",x"48",x"66",x"c4"),
  2386 => (x"7e",x"70",x"80",x"e0"),
  2387 => (x"c0",x"02",x"bf",x"6e"),
  2388 => (x"fd",x"4b",x"87",x"c5"),
  2389 => (x"c1",x"0f",x"73",x"49"),
  2390 => (x"49",x"fa",x"c3",x"7e"),
  2391 => (x"70",x"87",x"f8",x"e1"),
  2392 => (x"02",x"99",x"c2",x"49"),
  2393 => (x"c2",x"87",x"ea",x"c0"),
  2394 => (x"48",x"bf",x"c8",x"f7"),
  2395 => (x"03",x"a8",x"b7",x"c7"),
  2396 => (x"c2",x"87",x"c9",x"c0"),
  2397 => (x"c7",x"48",x"c8",x"f7"),
  2398 => (x"87",x"d3",x"c0",x"78"),
  2399 => (x"c1",x"48",x"66",x"c4"),
  2400 => (x"7e",x"70",x"80",x"e0"),
  2401 => (x"c0",x"02",x"bf",x"6e"),
  2402 => (x"fc",x"4b",x"87",x"c5"),
  2403 => (x"c1",x"0f",x"73",x"49"),
  2404 => (x"c3",x"48",x"75",x"7e"),
  2405 => (x"a6",x"cc",x"98",x"f0"),
  2406 => (x"05",x"98",x"70",x"58"),
  2407 => (x"c1",x"87",x"ce",x"c0"),
  2408 => (x"f2",x"e0",x"49",x"da"),
  2409 => (x"c2",x"49",x"70",x"87"),
  2410 => (x"f9",x"c1",x"02",x"99"),
  2411 => (x"49",x"e8",x"cf",x"87"),
  2412 => (x"70",x"87",x"cd",x"c3"),
  2413 => (x"c0",x"f7",x"c2",x"4b"),
  2414 => (x"c2",x"50",x"c0",x"48"),
  2415 => (x"bf",x"97",x"c0",x"f7"),
  2416 => (x"87",x"d2",x"c1",x"05"),
  2417 => (x"c0",x"05",x"66",x"c8"),
  2418 => (x"da",x"c1",x"87",x"cc"),
  2419 => (x"87",x"c7",x"e0",x"49"),
  2420 => (x"c1",x"02",x"98",x"70"),
  2421 => (x"bf",x"e8",x"87",x"c0"),
  2422 => (x"ff",x"c3",x"49",x"4d"),
  2423 => (x"2d",x"b7",x"c8",x"99"),
  2424 => (x"da",x"ff",x"b5",x"71"),
  2425 => (x"49",x"73",x"87",x"f4"),
  2426 => (x"70",x"87",x"e1",x"c2"),
  2427 => (x"c6",x"c0",x"02",x"98"),
  2428 => (x"c0",x"f7",x"c2",x"87"),
  2429 => (x"c2",x"50",x"c1",x"48"),
  2430 => (x"bf",x"97",x"c0",x"f7"),
  2431 => (x"87",x"d6",x"c0",x"05"),
  2432 => (x"f0",x"c3",x"49",x"75"),
  2433 => (x"cd",x"ff",x"05",x"99"),
  2434 => (x"49",x"da",x"c1",x"87"),
  2435 => (x"87",x"c7",x"df",x"ff"),
  2436 => (x"ff",x"05",x"98",x"70"),
  2437 => (x"f7",x"c2",x"87",x"c0"),
  2438 => (x"4b",x"49",x"bf",x"c8"),
  2439 => (x"66",x"c4",x"93",x"cc"),
  2440 => (x"71",x"4b",x"6b",x"83"),
  2441 => (x"9c",x"74",x"0f",x"73"),
  2442 => (x"87",x"e9",x"c0",x"02"),
  2443 => (x"e4",x"c0",x"02",x"6c"),
  2444 => (x"ff",x"49",x"6c",x"87"),
  2445 => (x"70",x"87",x"e0",x"de"),
  2446 => (x"02",x"99",x"c1",x"49"),
  2447 => (x"c4",x"87",x"cb",x"c0"),
  2448 => (x"f7",x"c2",x"4b",x"a4"),
  2449 => (x"6b",x"49",x"bf",x"c8"),
  2450 => (x"84",x"c8",x"0f",x"4b"),
  2451 => (x"87",x"c5",x"c0",x"02"),
  2452 => (x"dc",x"ff",x"05",x"6c"),
  2453 => (x"c0",x"02",x"6e",x"87"),
  2454 => (x"f7",x"c2",x"87",x"c8"),
  2455 => (x"f1",x"49",x"bf",x"c8"),
  2456 => (x"8e",x"f4",x"87",x"ea"),
  2457 => (x"4c",x"26",x"4d",x"26"),
  2458 => (x"4f",x"26",x"4b",x"26"),
  2459 => (x"00",x"00",x"00",x"10"),
  2460 => (x"00",x"00",x"00",x"00"),
  2461 => (x"00",x"00",x"00",x"00"),
  2462 => (x"00",x"00",x"00",x"00"),
  2463 => (x"00",x"00",x"00",x"00"),
  2464 => (x"ff",x"4a",x"71",x"1e"),
  2465 => (x"72",x"49",x"bf",x"c8"),
  2466 => (x"4f",x"26",x"48",x"a1"),
  2467 => (x"bf",x"c8",x"ff",x"1e"),
  2468 => (x"c0",x"c0",x"fe",x"89"),
  2469 => (x"a9",x"c0",x"c0",x"c0"),
  2470 => (x"c0",x"87",x"c4",x"01"),
  2471 => (x"c1",x"87",x"c2",x"4a"),
  2472 => (x"26",x"48",x"72",x"4a"),
  2473 => (x"5b",x"5e",x"0e",x"4f"),
  2474 => (x"71",x"0e",x"5d",x"5c"),
  2475 => (x"4c",x"d4",x"ff",x"4b"),
  2476 => (x"c0",x"48",x"66",x"d0"),
  2477 => (x"ff",x"49",x"d6",x"78"),
  2478 => (x"c3",x"87",x"d9",x"dd"),
  2479 => (x"49",x"6c",x"7c",x"ff"),
  2480 => (x"71",x"99",x"ff",x"c3"),
  2481 => (x"f0",x"c3",x"49",x"4d"),
  2482 => (x"a9",x"e0",x"c1",x"99"),
  2483 => (x"c3",x"87",x"cb",x"05"),
  2484 => (x"48",x"6c",x"7c",x"ff"),
  2485 => (x"66",x"d0",x"98",x"c3"),
  2486 => (x"ff",x"c3",x"78",x"08"),
  2487 => (x"49",x"4a",x"6c",x"7c"),
  2488 => (x"ff",x"c3",x"31",x"c8"),
  2489 => (x"71",x"4a",x"6c",x"7c"),
  2490 => (x"c8",x"49",x"72",x"b2"),
  2491 => (x"7c",x"ff",x"c3",x"31"),
  2492 => (x"b2",x"71",x"4a",x"6c"),
  2493 => (x"31",x"c8",x"49",x"72"),
  2494 => (x"6c",x"7c",x"ff",x"c3"),
  2495 => (x"ff",x"b2",x"71",x"4a"),
  2496 => (x"e0",x"c0",x"48",x"d0"),
  2497 => (x"02",x"9b",x"73",x"78"),
  2498 => (x"7b",x"72",x"87",x"c2"),
  2499 => (x"4d",x"26",x"48",x"75"),
  2500 => (x"4b",x"26",x"4c",x"26"),
  2501 => (x"26",x"1e",x"4f",x"26"),
  2502 => (x"5b",x"5e",x"0e",x"4f"),
  2503 => (x"86",x"f8",x"0e",x"5c"),
  2504 => (x"a6",x"c8",x"1e",x"76"),
  2505 => (x"87",x"fd",x"fd",x"49"),
  2506 => (x"4b",x"70",x"86",x"c4"),
  2507 => (x"a8",x"c4",x"48",x"6e"),
  2508 => (x"87",x"fb",x"c2",x"03"),
  2509 => (x"f0",x"c3",x"4a",x"73"),
  2510 => (x"aa",x"d0",x"c1",x"9a"),
  2511 => (x"c1",x"87",x"c7",x"02"),
  2512 => (x"c2",x"05",x"aa",x"e0"),
  2513 => (x"49",x"73",x"87",x"e9"),
  2514 => (x"c3",x"02",x"99",x"c8"),
  2515 => (x"87",x"c6",x"ff",x"87"),
  2516 => (x"9c",x"c3",x"4c",x"73"),
  2517 => (x"c1",x"05",x"ac",x"c2"),
  2518 => (x"66",x"c4",x"87",x"c4"),
  2519 => (x"71",x"31",x"c9",x"49"),
  2520 => (x"4a",x"66",x"c4",x"1e"),
  2521 => (x"c2",x"92",x"cc",x"c1"),
  2522 => (x"72",x"49",x"d0",x"f7"),
  2523 => (x"db",x"cd",x"fe",x"81"),
  2524 => (x"ff",x"49",x"d8",x"87"),
  2525 => (x"c8",x"87",x"dd",x"da"),
  2526 => (x"e4",x"c2",x"1e",x"c0"),
  2527 => (x"e6",x"fd",x"49",x"c8"),
  2528 => (x"d0",x"ff",x"87",x"f1"),
  2529 => (x"78",x"e0",x"c0",x"48"),
  2530 => (x"1e",x"c8",x"e4",x"c2"),
  2531 => (x"c1",x"4a",x"66",x"cc"),
  2532 => (x"f7",x"c2",x"92",x"cc"),
  2533 => (x"81",x"72",x"49",x"d0"),
  2534 => (x"87",x"f1",x"cb",x"fe"),
  2535 => (x"ac",x"c1",x"86",x"cc"),
  2536 => (x"87",x"cb",x"c1",x"05"),
  2537 => (x"fd",x"49",x"ee",x"c0"),
  2538 => (x"c4",x"87",x"e1",x"e3"),
  2539 => (x"31",x"c9",x"49",x"66"),
  2540 => (x"66",x"c4",x"1e",x"71"),
  2541 => (x"92",x"cc",x"c1",x"4a"),
  2542 => (x"49",x"d0",x"f7",x"c2"),
  2543 => (x"cc",x"fe",x"81",x"72"),
  2544 => (x"e4",x"c2",x"87",x"ca"),
  2545 => (x"66",x"c8",x"1e",x"c8"),
  2546 => (x"92",x"cc",x"c1",x"4a"),
  2547 => (x"49",x"d0",x"f7",x"c2"),
  2548 => (x"c9",x"fe",x"81",x"72"),
  2549 => (x"49",x"d7",x"87",x"f8"),
  2550 => (x"87",x"f8",x"d8",x"ff"),
  2551 => (x"c2",x"1e",x"c0",x"c8"),
  2552 => (x"fd",x"49",x"c8",x"e4"),
  2553 => (x"cc",x"87",x"e9",x"e4"),
  2554 => (x"48",x"d0",x"ff",x"86"),
  2555 => (x"f8",x"78",x"e0",x"c0"),
  2556 => (x"26",x"4c",x"26",x"8e"),
  2557 => (x"1e",x"4f",x"26",x"4b"),
  2558 => (x"b7",x"c4",x"4a",x"71"),
  2559 => (x"87",x"ce",x"03",x"aa"),
  2560 => (x"cc",x"c1",x"49",x"72"),
  2561 => (x"d0",x"f7",x"c2",x"91"),
  2562 => (x"81",x"c8",x"c1",x"81"),
  2563 => (x"4f",x"26",x"79",x"c0"),
  2564 => (x"5c",x"5b",x"5e",x"0e"),
  2565 => (x"86",x"fc",x"0e",x"5d"),
  2566 => (x"d4",x"ff",x"4a",x"71"),
  2567 => (x"d4",x"4c",x"c0",x"4b"),
  2568 => (x"b7",x"c3",x"4d",x"66"),
  2569 => (x"c2",x"c2",x"01",x"ad"),
  2570 => (x"02",x"9a",x"72",x"87"),
  2571 => (x"1e",x"87",x"ec",x"c0"),
  2572 => (x"cc",x"c1",x"49",x"75"),
  2573 => (x"d0",x"f7",x"c2",x"91"),
  2574 => (x"c8",x"80",x"71",x"48"),
  2575 => (x"66",x"c4",x"58",x"a6"),
  2576 => (x"d3",x"c3",x"fe",x"49"),
  2577 => (x"70",x"86",x"c4",x"87"),
  2578 => (x"87",x"d4",x"02",x"98"),
  2579 => (x"c8",x"c1",x"49",x"6e"),
  2580 => (x"6e",x"79",x"c1",x"81"),
  2581 => (x"69",x"81",x"c8",x"49"),
  2582 => (x"75",x"87",x"c5",x"4c"),
  2583 => (x"87",x"d7",x"fe",x"49"),
  2584 => (x"c8",x"48",x"d0",x"ff"),
  2585 => (x"7b",x"dd",x"78",x"e1"),
  2586 => (x"ff",x"c3",x"48",x"74"),
  2587 => (x"74",x"7b",x"70",x"98"),
  2588 => (x"29",x"b7",x"c8",x"49"),
  2589 => (x"ff",x"c3",x"48",x"71"),
  2590 => (x"74",x"7b",x"70",x"98"),
  2591 => (x"29",x"b7",x"d0",x"49"),
  2592 => (x"ff",x"c3",x"48",x"71"),
  2593 => (x"74",x"7b",x"70",x"98"),
  2594 => (x"28",x"b7",x"d8",x"48"),
  2595 => (x"7b",x"c0",x"7b",x"70"),
  2596 => (x"7b",x"7b",x"7b",x"7b"),
  2597 => (x"7b",x"7b",x"7b",x"7b"),
  2598 => (x"ff",x"7b",x"7b",x"7b"),
  2599 => (x"e0",x"c0",x"48",x"d0"),
  2600 => (x"dc",x"1e",x"75",x"78"),
  2601 => (x"d0",x"d6",x"ff",x"49"),
  2602 => (x"fc",x"86",x"c4",x"87"),
  2603 => (x"26",x"4d",x"26",x"8e"),
  2604 => (x"26",x"4b",x"26",x"4c"),
  2605 => (x"e3",x"c2",x"1e",x"4f"),
  2606 => (x"fe",x"49",x"bf",x"c4"),
  2607 => (x"c0",x"87",x"c3",x"dd"),
  2608 => (x"00",x"4f",x"26",x"48"),
  2609 => (x"00",x"00",x"28",x"c8"),
  2610 => (x"43",x"45",x"50",x"53"),
  2611 => (x"4d",x"55",x"52",x"54"),
  2612 => (x"00",x"4d",x"4f",x"52"),
  2613 => (x"00",x"00",x"1b",x"bf"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

